module hidden_layer_param (
    output reg signed [8*30*196-1:0] weights_HL, // Declare output as a flattened 1D array for weights
    output reg signed [8*30-1:0] biases_HL // Declare output as a flattened 1D array for biases
);

    // Local parameters for initialized weights and biases
    localparam signed [8*30*196-1:0] weights_HL_param = {
    8'sb00001011, 8'sb00001010, 8'sb00001011, 8'sb00001011, 8'sb00001100, 8'sb00001011, 8'sb00001110, 8'sb00001101, 8'sb00001011, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00001110, 8'sb00001100, 8'sb00001010, 8'sb00001010, 8'sb00001011, 8'sb00001101, 8'sb00010000, 8'sb00010001, 8'sb00010101, 8'sb00010010, 8'sb00010001, 8'sb00010001, 8'sb00010000, 8'sb00010001, 8'sb00001101, 8'sb00001010, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00001101, 8'sb00001001, 8'sb00010010, 8'sb00010111, 8'sb00011001, 8'sb00010111, 8'sb00011001, 8'sb00010100, 8'sb00001011, 8'sb00001101, 8'sb00001111, 8'sb00001110, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00001101, 8'sb00010000, 8'sb00010001, 8'sb00010101, 8'sb00001000, 8'sb00011000, 8'sb00010011, 8'sb00010000, 8'sb00010110, 8'sb00001101, 8'sb00001101, 8'sb00001100, 8'sb00001110, 8'sb00001111, 8'sb00001111, 8'sb00001011, 8'sb00001001, 8'sb00001101, 8'sb00010110, 8'sb00001111, 8'sb00011000, 8'sb00011010, 8'sb00100011, 8'sb00010010, 8'sb00001100, 8'sb00001110, 8'sb00001111, 8'sb00001000, 8'sb00000110, 8'sb00001101, 8'sb00001000, 8'sb00010011, 8'sb11111000, 8'sb11111111, 8'sb00001011, 8'sb00100000, 8'sb00100100, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00001010, 8'sb00001010, 8'sb00000010, 8'sb00011100, 8'sb00000100, 8'sb11110110, 8'sb11111111, 8'sb00000011, 8'sb00010111, 8'sb00010011, 8'sb00001011, 8'sb00001011, 8'sb00001110, 8'sb00000100, 8'sb00000011, 8'sb00001000, 8'sb00010000, 8'sb00011011, 8'sb00001010, 8'sb11111000, 8'sb11110001, 8'sb00000111, 8'sb00001010, 8'sb00001110, 8'sb00001001, 8'sb00001101, 8'sb00001110, 8'sb00000000, 8'sb11111100, 8'sb00001010, 8'sb00010100, 8'sb00011010, 8'sb11111010, 8'sb11110110, 8'sb11111100, 8'sb00001000, 8'sb00010011, 8'sb00001100, 8'sb00001010, 8'sb00001100, 8'sb00001101, 8'sb00001100, 8'sb00011100, 8'sb00010110, 8'sb00010010, 8'sb00001111, 8'sb11111100, 8'sb00010001, 8'sb00011010, 8'sb00010110, 8'sb00010101, 8'sb00001010, 8'sb00001010, 8'sb00001110, 8'sb00010000, 8'sb00011001, 8'sb00100111, 8'sb00100100, 8'sb00101010, 8'sb00110011, 8'sb00110010, 8'sb00101000, 8'sb00101111, 8'sb00101000, 8'sb00010101, 8'sb00000111, 8'sb00001011, 8'sb00001110, 8'sb00001110, 8'sb00010111, 8'sb00010100, 8'sb00011000, 8'sb00010111, 8'sb00100100, 8'sb00011110, 8'sb00100100, 8'sb00100110, 8'sb00100001, 8'sb00001101, 8'sb00001011, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00000110, 8'sb00001000, 8'sb00010101, 8'sb00010110, 8'sb00011101, 8'sb00011111, 8'sb00011100, 8'sb00010100, 8'sb00000111, 8'sb00001010, 8'sb00001100, 8'sb00001011, 8'sb00001010, 8'sb00001010, 8'sb00001100, 8'sb00001100, 8'sb00000111, 8'sb00001010, 8'sb00001011, 8'sb00001000, 8'sb00001100, 8'sb00001001, 8'sb00001100, 8'sb00001110, 8'sb00001101, 8'sb00001010,
    8'sb00001011, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001011, 8'sb00001100, 8'sb00001010, 8'sb00001011, 8'sb00001110, 8'sb00001010, 8'sb00001100, 8'sb00001101, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00001101, 8'sb00001010, 8'sb00001100, 8'sb00001001, 8'sb00001010, 8'sb00010010, 8'sb00001110, 8'sb00000110, 8'sb00000011, 8'sb00000111, 8'sb00000100, 8'sb00001010, 8'sb00001101, 8'sb00001100, 8'sb00001101, 8'sb00001100, 8'sb00010000, 8'sb00010100, 8'sb00011010, 8'sb00011001, 8'sb00011010, 8'sb00100100, 8'sb00011111, 8'sb00001010, 8'sb00000001, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001100, 8'sb00010100, 8'sb00011000, 8'sb00001111, 8'sb00010001, 8'sb00010101, 8'sb00001100, 8'sb00001011, 8'sb00011111, 8'sb00011011, 8'sb00011000, 8'sb00010110, 8'sb00001101, 8'sb00001101, 8'sb00001010, 8'sb00010010, 8'sb00010010, 8'sb00010010, 8'sb00100010, 8'sb00100000, 8'sb00010011, 8'sb00010010, 8'sb00011010, 8'sb00011001, 8'sb00100010, 8'sb00100011, 8'sb00010010, 8'sb00001101, 8'sb00001100, 8'sb00001110, 8'sb00001011, 8'sb00000100, 8'sb00000111, 8'sb00010001, 8'sb00010001, 8'sb00000000, 8'sb00001110, 8'sb00001110, 8'sb00010011, 8'sb00100000, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00000110, 8'sb00000101, 8'sb00000100, 8'sb11111110, 8'sb00011110, 8'sb00010000, 8'sb00000011, 8'sb00001101, 8'sb11111100, 8'sb11110100, 8'sb00000010, 8'sb00001101, 8'sb00001010, 8'sb00001100, 8'sb00001011, 8'sb00000111, 8'sb00001110, 8'sb00000011, 8'sb00010101, 8'sb00001000, 8'sb11111100, 8'sb11111101, 8'sb11111010, 8'sb00000010, 8'sb00001001, 8'sb00010000, 8'sb00001100, 8'sb00010000, 8'sb00010101, 8'sb11111110, 8'sb00000100, 8'sb00001010, 8'sb00001110, 8'sb00000000, 8'sb00000101, 8'sb00001010, 8'sb00010011, 8'sb00011011, 8'sb00010100, 8'sb00001100, 8'sb00001100, 8'sb00001111, 8'sb00011110, 8'sb00010001, 8'sb00010000, 8'sb00010001, 8'sb00000000, 8'sb00011001, 8'sb00011011, 8'sb00011010, 8'sb00011010, 8'sb00100111, 8'sb00010111, 8'sb00001110, 8'sb00001011, 8'sb00001111, 8'sb00011011, 8'sb00100101, 8'sb00010011, 8'sb00010000, 8'sb00000101, 8'sb00010000, 8'sb00010011, 8'sb00010001, 8'sb00100001, 8'sb00100001, 8'sb00010000, 8'sb00001100, 8'sb00001010, 8'sb00010000, 8'sb00010100, 8'sb00011101, 8'sb00001101, 8'sb00010000, 8'sb00001110, 8'sb00000111, 8'sb00010101, 8'sb00010001, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00001101, 8'sb00001010, 8'sb00001110, 8'sb00001001, 8'sb00000101, 8'sb00010010, 8'sb00010100, 8'sb00011000, 8'sb00010101, 8'sb00010110, 8'sb00001110, 8'sb00000101, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00001011, 8'sb00001100, 8'sb00001100, 8'sb00001101, 8'sb00010000, 8'sb00010010, 8'sb00010011, 8'sb00001011, 8'sb00001001, 8'sb00001100, 8'sb00001100, 8'sb00001101,
    8'sb00010001, 8'sb00001101, 8'sb00001111, 8'sb00010001, 8'sb00001101, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00001111, 8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00001100, 8'sb00001100, 8'sb00010001, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010011, 8'sb00010101, 8'sb00011010, 8'sb00010101, 8'sb00010111, 8'sb00010011, 8'sb00001110, 8'sb00001100, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00010001, 8'sb00010100, 8'sb00011101, 8'sb00100100, 8'sb00011010, 8'sb00010011, 8'sb00010011, 8'sb00010100, 8'sb00010101, 8'sb00001010, 8'sb00001010, 8'sb00001101, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00011100, 8'sb00100100, 8'sb00010111, 8'sb00001111, 8'sb00010111, 8'sb00001011, 8'sb00001110, 8'sb00001111, 8'sb00001001, 8'sb00000100, 8'sb00000010, 8'sb00001101, 8'sb00010000, 8'sb00010010, 8'sb00100000, 8'sb00001000, 8'sb00000000, 8'sb00000000, 8'sb00001000, 8'sb00010111, 8'sb00100001, 8'sb00001110, 8'sb00001101, 8'sb00000100, 8'sb11110111, 8'sb00001001, 8'sb00001100, 8'sb00010010, 8'sb00000110, 8'sb11100010, 8'sb11101101, 8'sb11110001, 8'sb11111011, 8'sb11110110, 8'sb00011011, 8'sb00010011, 8'sb00010110, 8'sb00010000, 8'sb00000011, 8'sb00001011, 8'sb00010000, 8'sb00001110, 8'sb11111111, 8'sb00000100, 8'sb00001111, 8'sb00001100, 8'sb00001111, 8'sb11110110, 8'sb00010010, 8'sb11111110, 8'sb00000000, 8'sb00100100, 8'sb00100010, 8'sb00001110, 8'sb00001110, 8'sb00001111, 8'sb00011001, 8'sb00100000, 8'sb00011001, 8'sb00010001, 8'sb00000111, 8'sb11110101, 8'sb00010000, 8'sb00001010, 8'sb00011000, 8'sb00100011, 8'sb00011010, 8'sb00001111, 8'sb00001100, 8'sb00010001, 8'sb00010001, 8'sb00011100, 8'sb00011101, 8'sb00010000, 8'sb00001001, 8'sb00001000, 8'sb00011110, 8'sb00011111, 8'sb00011110, 8'sb00100000, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00010110, 8'sb00001101, 8'sb00010000, 8'sb00010000, 8'sb00010010, 8'sb00001000, 8'sb00010111, 8'sb00011110, 8'sb00011010, 8'sb00011001, 8'sb00010010, 8'sb00001100, 8'sb00010001, 8'sb00010000, 8'sb00010101, 8'sb00010011, 8'sb00010111, 8'sb00010001, 8'sb00010110, 8'sb00010111, 8'sb00010010, 8'sb00010100, 8'sb00010110, 8'sb00010101, 8'sb00000011, 8'sb00001101, 8'sb00001111, 8'sb00001101, 8'sb00010011, 8'sb00010000, 8'sb00010010, 8'sb00010000, 8'sb00010101, 8'sb00001111, 8'sb00010001, 8'sb00000111, 8'sb00001010, 8'sb00000101, 8'sb00001001, 8'sb00001101, 8'sb00001100, 8'sb00001110, 8'sb00010000, 8'sb00010110, 8'sb00011001, 8'sb00011001, 8'sb00010110, 8'sb00010011, 8'sb00001110, 8'sb00001111, 8'sb00000000, 8'sb00000010, 8'sb00001011, 8'sb00010000, 8'sb00010001, 8'sb00001100, 8'sb00010001, 8'sb00001101, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00010000, 8'sb00001101, 8'sb00010000, 8'sb00001111, 8'sb00001110, 8'sb00001111, 8'sb00001110,
    8'sb00001111, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00010011, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010011, 8'sb00001111, 8'sb00001111, 8'sb00010000, 8'sb00001101, 8'sb00001110, 8'sb00001111, 8'sb00010001, 8'sb00010010, 8'sb00001111, 8'sb00010010, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00010100, 8'sb00010001, 8'sb00001101, 8'sb00010110, 8'sb00010000, 8'sb00001101, 8'sb00001111, 8'sb00001101, 8'sb00010000, 8'sb00011000, 8'sb00010110, 8'sb00010010, 8'sb00010010, 8'sb00010010, 8'sb00010111, 8'sb00001101, 8'sb00010100, 8'sb00010010, 8'sb00010100, 8'sb00010010, 8'sb00010101, 8'sb00010010, 8'sb00010100, 8'sb00010010, 8'sb00011110, 8'sb00010101, 8'sb00010010, 8'sb00010101, 8'sb00010100, 8'sb00010000, 8'sb00011001, 8'sb00010011, 8'sb00010011, 8'sb00001110, 8'sb00001101, 8'sb00001010, 8'sb00001011, 8'sb00001101, 8'sb00011101, 8'sb00010100, 8'sb00010011, 8'sb00010110, 8'sb00001101, 8'sb00000111, 8'sb00000110, 8'sb00000100, 8'sb00001101, 8'sb11111111, 8'sb00000010, 8'sb00000110, 8'sb00000000, 8'sb11111011, 8'sb00001011, 8'sb00010001, 8'sb00010011, 8'sb00010110, 8'sb00010001, 8'sb00001001, 8'sb00010000, 8'sb00001111, 8'sb00010110, 8'sb00001110, 8'sb00010000, 8'sb00001100, 8'sb00000100, 8'sb11111100, 8'sb00000011, 8'sb00001111, 8'sb00010000, 8'sb00010000, 8'sb00001101, 8'sb00000110, 8'sb00011000, 8'sb00010110, 8'sb00010111, 8'sb00010001, 8'sb00000101, 8'sb00001001, 8'sb00010000, 8'sb00011000, 8'sb00001110, 8'sb00010000, 8'sb00010011, 8'sb00010100, 8'sb11111010, 8'sb11011011, 8'sb11101000, 8'sb00001010, 8'sb00011100, 8'sb00000100, 8'sb00001010, 8'sb00011000, 8'sb00010010, 8'sb00011010, 8'sb00010100, 8'sb00010001, 8'sb00010010, 8'sb00011001, 8'sb00000001, 8'sb11101110, 8'sb11011100, 8'sb11000010, 8'sb11001001, 8'sb11111011, 8'sb00001110, 8'sb00010001, 8'sb00010001, 8'sb00010011, 8'sb00010001, 8'sb00010001, 8'sb00010010, 8'sb00010111, 8'sb00010110, 8'sb00001110, 8'sb00010111, 8'sb00100001, 8'sb00100000, 8'sb00010100, 8'sb00001000, 8'sb00001011, 8'sb00010000, 8'sb00001100, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00010010, 8'sb00011100, 8'sb00011011, 8'sb00010111, 8'sb00011110, 8'sb00011100, 8'sb00011100, 8'sb00010011, 8'sb00010010, 8'sb00001001, 8'sb00001111, 8'sb00001111, 8'sb00010010, 8'sb00010000, 8'sb00010001, 8'sb00011000, 8'sb00101001, 8'sb00100101, 8'sb00011110, 8'sb00011000, 8'sb00010011, 8'sb00010001, 8'sb00001011, 8'sb00010000, 8'sb00010101, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00010001, 8'sb00010000, 8'sb00010100, 8'sb00010001, 8'sb00010110, 8'sb00010100, 8'sb00010010, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00010011,
    8'sb00001010, 8'sb00001100, 8'sb00001011, 8'sb00001011, 8'sb00001011, 8'sb00001100, 8'sb00001100, 8'sb00001101, 8'sb00001110, 8'sb00001011, 8'sb00001011, 8'sb00001100, 8'sb00001111, 8'sb00001100, 8'sb00001010, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00001011, 8'sb00001011, 8'sb00001011, 8'sb00001101, 8'sb00001101, 8'sb00010001, 8'sb00010001, 8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00001011, 8'sb00001011, 8'sb00001111, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00001001, 8'sb00000100, 8'sb00001000, 8'sb00010011, 8'sb00010001, 8'sb00010001, 8'sb00010000, 8'sb00001101, 8'sb00001100, 8'sb00001011, 8'sb00010011, 8'sb00010011, 8'sb00010101, 8'sb00010011, 8'sb00010000, 8'sb00001101, 8'sb00001111, 8'sb00011101, 8'sb00001111, 8'sb00001110, 8'sb00010010, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00010000, 8'sb00010010, 8'sb00001011, 8'sb00001110, 8'sb00001001, 8'sb00001011, 8'sb00001100, 8'sb00001110, 8'sb00011100, 8'sb00011001, 8'sb00011001, 8'sb00001111, 8'sb00001010, 8'sb00001100, 8'sb00010000, 8'sb00010001, 8'sb00001001, 8'sb00001101, 8'sb00001110, 8'sb00001101, 8'sb00100000, 8'sb00000100, 8'sb11111101, 8'sb00000010, 8'sb00001000, 8'sb00001110, 8'sb00001100, 8'sb00001111, 8'sb00011011, 8'sb00010111, 8'sb00010011, 8'sb00010110, 8'sb00001101, 8'sb00010100, 8'sb00100101, 8'sb00011100, 8'sb00001010, 8'sb11111000, 8'sb11111110, 8'sb00001010, 8'sb00001110, 8'sb00001110, 8'sb00001111, 8'sb00000100, 8'sb11111001, 8'sb11111110, 8'sb00000100, 8'sb00011011, 8'sb00011011, 8'sb00011000, 8'sb00011101, 8'sb00010000, 8'sb00000101, 8'sb00001011, 8'sb00001100, 8'sb00001111, 8'sb00000101, 8'sb00000101, 8'sb00000000, 8'sb11100110, 8'sb00001111, 8'sb00100001, 8'sb00001110, 8'sb00011001, 8'sb00010100, 8'sb00000110, 8'sb00000100, 8'sb00001011, 8'sb00001100, 8'sb00010011, 8'sb00001111, 8'sb00001111, 8'sb00000010, 8'sb11101011, 8'sb00100001, 8'sb00011101, 8'sb00011000, 8'sb00010111, 8'sb00010000, 8'sb11111110, 8'sb00000001, 8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00001101, 8'sb00000010, 8'sb11111101, 8'sb11111100, 8'sb00001111, 8'sb00011010, 8'sb00101001, 8'sb00010110, 8'sb00001111, 8'sb00001001, 8'sb00001010, 8'sb00001011, 8'sb00001100, 8'sb00001011, 8'sb00001111, 8'sb11111100, 8'sb11111110, 8'sb00000110, 8'sb11111101, 8'sb00001111, 8'sb00010111, 8'sb00010110, 8'sb00010010, 8'sb00010001, 8'sb00001111, 8'sb00001101, 8'sb00001011, 8'sb00001110, 8'sb00010111, 8'sb00100010, 8'sb00011000, 8'sb00001100, 8'sb00001010, 8'sb00010010, 8'sb00010110, 8'sb00010111, 8'sb00010111, 8'sb00010011, 8'sb00001010, 8'sb00001100, 8'sb00001011, 8'sb00001110, 8'sb00001101, 8'sb00010000, 8'sb00010010, 8'sb00010000, 8'sb00010010, 8'sb00010001, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001100, 8'sb00001101,
    8'sb00010100, 8'sb00010011, 8'sb00010011, 8'sb00010011, 8'sb00010000, 8'sb00010001, 8'sb00010000, 8'sb00010100, 8'sb00010000, 8'sb00010000, 8'sb00010011, 8'sb00010100, 8'sb00010000, 8'sb00010100, 8'sb00010010, 8'sb00010011, 8'sb00010001, 8'sb00010011, 8'sb00010111, 8'sb00011010, 8'sb00011000, 8'sb00010001, 8'sb00010000, 8'sb00001101, 8'sb00001011, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00010100, 8'sb00010011, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00011000, 8'sb00001100, 8'sb00001010, 8'sb00001000, 8'sb00010000, 8'sb00010100, 8'sb00010100, 8'sb00010010, 8'sb00001101, 8'sb00000001, 8'sb00000110, 8'sb00001110, 8'sb00000111, 8'sb00010100, 8'sb00010100, 8'sb00010000, 8'sb00010001, 8'sb00001010, 8'sb00000100, 8'sb00010010, 8'sb00010001, 8'sb00010000, 8'sb00001101, 8'sb00001010, 8'sb00010001, 8'sb00011001, 8'sb00000110, 8'sb00001001, 8'sb00010000, 8'sb00001001, 8'sb00001000, 8'sb11111101, 8'sb11111101, 8'sb00010100, 8'sb00010001, 8'sb00010000, 8'sb00001001, 8'sb11111110, 8'sb00000110, 8'sb11111110, 8'sb11110100, 8'sb00000110, 8'sb00011010, 8'sb00000110, 8'sb00001100, 8'sb11111100, 8'sb00001101, 8'sb00010010, 8'sb00010011, 8'sb00010010, 8'sb11110111, 8'sb11011111, 8'sb11100101, 8'sb11110011, 8'sb00000001, 8'sb00000001, 8'sb00000111, 8'sb00000111, 8'sb00010000, 8'sb00000000, 8'sb00001110, 8'sb00010101, 8'sb00010010, 8'sb00010100, 8'sb00000101, 8'sb00001101, 8'sb00011100, 8'sb00011110, 8'sb00011101, 8'sb00001010, 8'sb00000101, 8'sb11110110, 8'sb11110110, 8'sb00000100, 8'sb00011000, 8'sb00011000, 8'sb00010001, 8'sb00010011, 8'sb00011100, 8'sb00011101, 8'sb00010111, 8'sb00010110, 8'sb00101010, 8'sb00010000, 8'sb11111110, 8'sb00000000, 8'sb00010010, 8'sb00011011, 8'sb00100110, 8'sb00010111, 8'sb00010010, 8'sb00001111, 8'sb00011001, 8'sb00010110, 8'sb00011101, 8'sb00011101, 8'sb00101001, 8'sb11110001, 8'sb00000001, 8'sb00001100, 8'sb00010110, 8'sb00011001, 8'sb00100111, 8'sb00010110, 8'sb00010001, 8'sb00010010, 8'sb00011011, 8'sb00010000, 8'sb00010110, 8'sb00011000, 8'sb00000111, 8'sb00000000, 8'sb00001010, 8'sb00010110, 8'sb00001000, 8'sb00010111, 8'sb00011100, 8'sb00010011, 8'sb00010010, 8'sb00010001, 8'sb00011010, 8'sb00001110, 8'sb00001100, 8'sb00001000, 8'sb00001111, 8'sb00000110, 8'sb00001010, 8'sb00011010, 8'sb00010110, 8'sb00010101, 8'sb00010011, 8'sb00010011, 8'sb00010100, 8'sb00010001, 8'sb00001101, 8'sb00000010, 8'sb11111110, 8'sb00000011, 8'sb00001110, 8'sb00001101, 8'sb00001011, 8'sb00001001, 8'sb00010000, 8'sb00010001, 8'sb00010100, 8'sb00010101, 8'sb00010100, 8'sb00010011, 8'sb00010101, 8'sb00001111, 8'sb00010001, 8'sb00010001, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00010100, 8'sb00010001, 8'sb00010010,
    8'sb00010100, 8'sb00010010, 8'sb00010011, 8'sb00010000, 8'sb00010100, 8'sb00010000, 8'sb00010010, 8'sb00010000, 8'sb00010000, 8'sb00010100, 8'sb00010001, 8'sb00010010, 8'sb00010011, 8'sb00010101, 8'sb00010100, 8'sb00010100, 8'sb00010010, 8'sb00010000, 8'sb00001111, 8'sb00001010, 8'sb00000111, 8'sb00000010, 8'sb00000101, 8'sb00001101, 8'sb00001100, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00010101, 8'sb00010001, 8'sb00000111, 8'sb11111110, 8'sb11111011, 8'sb11111101, 8'sb00000000, 8'sb11111001, 8'sb11111010, 8'sb00000001, 8'sb00001010, 8'sb00001110, 8'sb00010011, 8'sb00010101, 8'sb00010011, 8'sb00010101, 8'sb00001011, 8'sb00001001, 8'sb00001000, 8'sb00000011, 8'sb00001110, 8'sb00010001, 8'sb00001110, 8'sb00010101, 8'sb00011010, 8'sb00011100, 8'sb00010011, 8'sb00010010, 8'sb00011001, 8'sb00010110, 8'sb00010001, 8'sb00010001, 8'sb11111011, 8'sb00010101, 8'sb00010101, 8'sb00100001, 8'sb00011100, 8'sb00010111, 8'sb00011010, 8'sb00100000, 8'sb00010110, 8'sb00010001, 8'sb00010111, 8'sb00001100, 8'sb00000001, 8'sb00001110, 8'sb00100000, 8'sb00010010, 8'sb00010100, 8'sb00010110, 8'sb00001101, 8'sb00010001, 8'sb00011110, 8'sb00100011, 8'sb00010110, 8'sb00010101, 8'sb00010110, 8'sb00010010, 8'sb00011111, 8'sb00100001, 8'sb00011001, 8'sb00000001, 8'sb00010010, 8'sb00010000, 8'sb00000010, 8'sb11111110, 8'sb11111100, 8'sb00001011, 8'sb00010011, 8'sb00010010, 8'sb00010110, 8'sb00010000, 8'sb00010001, 8'sb00010110, 8'sb00000110, 8'sb00001000, 8'sb00010000, 8'sb00100101, 8'sb00001110, 8'sb00001110, 8'sb00000111, 8'sb00001010, 8'sb00010011, 8'sb00010001, 8'sb00001101, 8'sb11111111, 8'sb00000101, 8'sb00010100, 8'sb00010010, 8'sb00010111, 8'sb00010101, 8'sb00001011, 8'sb00000110, 8'sb00001100, 8'sb11111100, 8'sb00000001, 8'sb00001111, 8'sb00010011, 8'sb00001110, 8'sb11110010, 8'sb11111011, 8'sb00000110, 8'sb00001101, 8'sb00011011, 8'sb00001110, 8'sb11111011, 8'sb00000101, 8'sb00000001, 8'sb11110000, 8'sb00000010, 8'sb00010011, 8'sb00010010, 8'sb00001110, 8'sb11110100, 8'sb11111100, 8'sb00000010, 8'sb11111100, 8'sb00000100, 8'sb00001011, 8'sb00000010, 8'sb11111110, 8'sb11111111, 8'sb00000101, 8'sb00001100, 8'sb00010001, 8'sb00010001, 8'sb00001111, 8'sb00001101, 8'sb00001110, 8'sb00001111, 8'sb00010000, 8'sb00001010, 8'sb00001100, 8'sb00001000, 8'sb00000100, 8'sb00000001, 8'sb00010001, 8'sb00010010, 8'sb00010100, 8'sb00010100, 8'sb00010101, 8'sb00010001, 8'sb00010101, 8'sb00010001, 8'sb00001101, 8'sb00001010, 8'sb00010001, 8'sb00001010, 8'sb00010010, 8'sb00010001, 8'sb00010101, 8'sb00010000, 8'sb00010100, 8'sb00010001, 8'sb00010001, 8'sb00010101, 8'sb00010100, 8'sb00010011, 8'sb00010100, 8'sb00010100, 8'sb00010111, 8'sb00010001, 8'sb00010011, 8'sb00010001, 8'sb00010100, 8'sb00010001, 8'sb00010010,
    8'sb00001111, 8'sb00010001, 8'sb00010001, 8'sb00010011, 8'sb00010001, 8'sb00010100, 8'sb00010100, 8'sb00010011, 8'sb00010001, 8'sb00010000, 8'sb00010000, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00010001, 8'sb00010001, 8'sb00010010, 8'sb00010001, 8'sb00011000, 8'sb00010110, 8'sb00010101, 8'sb00011010, 8'sb00010011, 8'sb00010001, 8'sb00001101, 8'sb00010000, 8'sb00010001, 8'sb00010011, 8'sb00010011, 8'sb00010011, 8'sb00010000, 8'sb00010010, 8'sb00001111, 8'sb00001110, 8'sb00011000, 8'sb00011000, 8'sb00000101, 8'sb00000011, 8'sb00001010, 8'sb00001101, 8'sb00001111, 8'sb00010001, 8'sb00010010, 8'sb00010011, 8'sb00010000, 8'sb00011001, 8'sb00001101, 8'sb00001110, 8'sb00000101, 8'sb11110100, 8'sb00001001, 8'sb00001010, 8'sb00000111, 8'sb00000100, 8'sb00001010, 8'sb00001110, 8'sb00010100, 8'sb00011010, 8'sb00011001, 8'sb00010111, 8'sb00001111, 8'sb00010010, 8'sb00001011, 8'sb00001010, 8'sb00001000, 8'sb00001100, 8'sb00001011, 8'sb00001110, 8'sb00000111, 8'sb00001111, 8'sb00010010, 8'sb00011100, 8'sb00011011, 8'sb00010010, 8'sb00010010, 8'sb00011011, 8'sb00001101, 8'sb00001000, 8'sb00001101, 8'sb00001101, 8'sb00010010, 8'sb00010000, 8'sb00001101, 8'sb00001110, 8'sb00010010, 8'sb00011011, 8'sb00011010, 8'sb00011001, 8'sb00011101, 8'sb00001011, 8'sb11100011, 8'sb00001010, 8'sb00000110, 8'sb00010000, 8'sb00001100, 8'sb00010011, 8'sb00010101, 8'sb00010000, 8'sb00010000, 8'sb00010011, 8'sb00001011, 8'sb00001110, 8'sb00000101, 8'sb11011111, 8'sb00000001, 8'sb00010101, 8'sb00000110, 8'sb00001101, 8'sb00001110, 8'sb00011101, 8'sb00010110, 8'sb00010000, 8'sb00001111, 8'sb00001110, 8'sb00000110, 8'sb00000010, 8'sb11100101, 8'sb11011101, 8'sb00100010, 8'sb00011110, 8'sb00010101, 8'sb00001110, 8'sb00010010, 8'sb00001110, 8'sb00011000, 8'sb00010000, 8'sb00010011, 8'sb00010000, 8'sb00000100, 8'sb11110101, 8'sb11101010, 8'sb11111101, 8'sb00111011, 8'sb00011110, 8'sb00010100, 8'sb00010100, 8'sb00000110, 8'sb00001000, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00010000, 8'sb00000010, 8'sb11111101, 8'sb11111100, 8'sb00010110, 8'sb00100100, 8'sb00100100, 8'sb00010111, 8'sb00010101, 8'sb00000010, 8'sb00001010, 8'sb00010010, 8'sb00010100, 8'sb00010000, 8'sb00010001, 8'sb00001101, 8'sb00001010, 8'sb00000110, 8'sb11111100, 8'sb00001000, 8'sb00010000, 8'sb00011011, 8'sb00011001, 8'sb00001000, 8'sb00001001, 8'sb00010010, 8'sb00010010, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00001011, 8'sb00001010, 8'sb00000101, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00001100, 8'sb00001101, 8'sb00010001, 8'sb00001111, 8'sb00010011, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00010100, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00010010, 8'sb00011001, 8'sb00010100, 8'sb00010011, 8'sb00010001, 8'sb00010001,
    8'sb00001111, 8'sb00001101, 8'sb00001101, 8'sb00001011, 8'sb00001011, 8'sb00001100, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00001011, 8'sb00010000, 8'sb00001100, 8'sb00001110, 8'sb00001111, 8'sb00001110, 8'sb00000111, 8'sb11111111, 8'sb00000010, 8'sb11111110, 8'sb00001001, 8'sb00010100, 8'sb00001111, 8'sb00001011, 8'sb00001011, 8'sb00001100, 8'sb00001110, 8'sb00010000, 8'sb00010000, 8'sb00010001, 8'sb00001011, 8'sb00001100, 8'sb00001101, 8'sb00010011, 8'sb00000011, 8'sb11111111, 8'sb00000001, 8'sb00010010, 8'sb00011001, 8'sb00010101, 8'sb00010001, 8'sb00001100, 8'sb00001101, 8'sb00010110, 8'sb00010100, 8'sb00011000, 8'sb00011001, 8'sb00010111, 8'sb00011011, 8'sb00011101, 8'sb00011100, 8'sb00011101, 8'sb00101001, 8'sb00010101, 8'sb00001101, 8'sb00001111, 8'sb00010010, 8'sb00010000, 8'sb00010001, 8'sb00010100, 8'sb00010000, 8'sb00011101, 8'sb00011111, 8'sb00110000, 8'sb00100101, 8'sb00011010, 8'sb00011100, 8'sb00001101, 8'sb00001010, 8'sb00001111, 8'sb00010001, 8'sb00001110, 8'sb00010011, 8'sb00010111, 8'sb00011001, 8'sb00010101, 8'sb00001000, 8'sb00001111, 8'sb00001100, 8'sb00011000, 8'sb00010010, 8'sb00001101, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00011001, 8'sb00101011, 8'sb00100111, 8'sb00100010, 8'sb00010100, 8'sb00000011, 8'sb00001011, 8'sb00010010, 8'sb00001110, 8'sb00010110, 8'sb00001110, 8'sb00001111, 8'sb00001111, 8'sb00001100, 8'sb00011110, 8'sb00010110, 8'sb00011000, 8'sb00010100, 8'sb00000101, 8'sb00000111, 8'sb00010000, 8'sb00010010, 8'sb00001000, 8'sb00001110, 8'sb00001000, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00000011, 8'sb00001000, 8'sb00010111, 8'sb00010000, 8'sb00010010, 8'sb00000101, 8'sb00010110, 8'sb00010001, 8'sb00001110, 8'sb00010010, 8'sb00000010, 8'sb00001101, 8'sb00010000, 8'sb00001011, 8'sb11111110, 8'sb00000110, 8'sb11111111, 8'sb00000000, 8'sb11111111, 8'sb11111101, 8'sb00001010, 8'sb00001101, 8'sb00001000, 8'sb00001000, 8'sb11111110, 8'sb00001111, 8'sb00001111, 8'sb00001101, 8'sb00000000, 8'sb11111101, 8'sb11111000, 8'sb11110111, 8'sb11111101, 8'sb11111111, 8'sb00000111, 8'sb00000010, 8'sb00010000, 8'sb00000000, 8'sb00000100, 8'sb00001011, 8'sb00001110, 8'sb00001110, 8'sb00001001, 8'sb00010101, 8'sb00001111, 8'sb00010011, 8'sb00011010, 8'sb00010100, 8'sb00010001, 8'sb00001010, 8'sb00010001, 8'sb00001001, 8'sb00001011, 8'sb00001111, 8'sb00001110, 8'sb00001111, 8'sb00010011, 8'sb00011011, 8'sb00011110, 8'sb00100101, 8'sb00100100, 8'sb00100101, 8'sb00011101, 8'sb00010001, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00001100, 8'sb00010000, 8'sb00001101, 8'sb00010000, 8'sb00010010, 8'sb00010011, 8'sb00001101, 8'sb00001111, 8'sb00001111, 8'sb00010000, 8'sb00001110, 8'sb00001111,
    8'sb00010000, 8'sb00010010, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00010010, 8'sb00001111, 8'sb00001110, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010110, 8'sb00011111, 8'sb00011100, 8'sb00010010, 8'sb00000100, 8'sb00000101, 8'sb00000111, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00001110, 8'sb00010001, 8'sb00011000, 8'sb00011001, 8'sb00100000, 8'sb00100100, 8'sb00011110, 8'sb00001110, 8'sb00001100, 8'sb00000000, 8'sb00000001, 8'sb00010010, 8'sb00001111, 8'sb00001111, 8'sb00001111, 8'sb00010011, 8'sb00001001, 8'sb00000101, 8'sb00010011, 8'sb00100100, 8'sb00011111, 8'sb00011011, 8'sb00001100, 8'sb00011100, 8'sb00010110, 8'sb00010110, 8'sb00010011, 8'sb00010010, 8'sb00001111, 8'sb00010000, 8'sb00001100, 8'sb00000111, 8'sb00000000, 8'sb00011011, 8'sb00101001, 8'sb00010111, 8'sb00010001, 8'sb00011010, 8'sb00011101, 8'sb00010110, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00001111, 8'sb11111111, 8'sb11111001, 8'sb11100101, 8'sb11101111, 8'sb00011111, 8'sb00011000, 8'sb00010100, 8'sb00000101, 8'sb00000011, 8'sb00010100, 8'sb00001110, 8'sb00001101, 8'sb00001110, 8'sb11111001, 8'sb11100010, 8'sb11111010, 8'sb11111101, 8'sb11111001, 8'sb00011000, 8'sb00000101, 8'sb00001011, 8'sb00000101, 8'sb11111001, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00001111, 8'sb00001010, 8'sb00001010, 8'sb00010000, 8'sb00001010, 8'sb00010001, 8'sb00011011, 8'sb00001010, 8'sb00001100, 8'sb00000100, 8'sb00000010, 8'sb00010101, 8'sb00010100, 8'sb00010001, 8'sb00010110, 8'sb00100010, 8'sb00001010, 8'sb00000100, 8'sb11111100, 8'sb00000001, 8'sb00010000, 8'sb00000101, 8'sb00001001, 8'sb00000111, 8'sb00000111, 8'sb00011000, 8'sb00010001, 8'sb00010001, 8'sb00010100, 8'sb00101001, 8'sb00011001, 8'sb00010111, 8'sb00000101, 8'sb00001110, 8'sb00010111, 8'sb00010010, 8'sb00011001, 8'sb00010001, 8'sb00010111, 8'sb00100000, 8'sb00001111, 8'sb00010000, 8'sb00010100, 8'sb00100001, 8'sb00100101, 8'sb00011101, 8'sb00011001, 8'sb00010000, 8'sb00010001, 8'sb00010100, 8'sb00010110, 8'sb00011000, 8'sb00011001, 8'sb00010110, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00010001, 8'sb00010110, 8'sb00011000, 8'sb00010111, 8'sb00000100, 8'sb00001000, 8'sb00001100, 8'sb00010100, 8'sb00010001, 8'sb00010101, 8'sb00010100, 8'sb00010010, 8'sb00001111, 8'sb00010011, 8'sb00010001, 8'sb00001100, 8'sb00001100, 8'sb00001101, 8'sb00010110, 8'sb00001100, 8'sb00001000, 8'sb00000100, 8'sb00000110, 8'sb00001110, 8'sb00010011, 8'sb00010000, 8'sb00001110, 8'sb00001111, 8'sb00001110, 8'sb00010000, 8'sb00001101, 8'sb00001101, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00010001, 8'sb00001110, 8'sb00001110, 8'sb00010001, 8'sb00001110,
    8'sb00010000, 8'sb00001111, 8'sb00001101, 8'sb00001101, 8'sb00001101, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00001011, 8'sb00001011, 8'sb00001010, 8'sb00001011, 8'sb00001110, 8'sb00011000, 8'sb00010111, 8'sb00010010, 8'sb00001101, 8'sb00010000, 8'sb00001101, 8'sb00001110, 8'sb00010000, 8'sb00001111, 8'sb00001001, 8'sb00001101, 8'sb00001001, 8'sb00001101, 8'sb00010100, 8'sb00100101, 8'sb00100011, 8'sb00100000, 8'sb00011011, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00001011, 8'sb00001100, 8'sb00010001, 8'sb00011001, 8'sb11111001, 8'sb11110001, 8'sb11110111, 8'sb11111100, 8'sb00000011, 8'sb00000110, 8'sb00101001, 8'sb00011000, 8'sb00001111, 8'sb00010000, 8'sb00001011, 8'sb00000111, 8'sb00000100, 8'sb00000110, 8'sb11111011, 8'sb11101011, 8'sb11101101, 8'sb00000100, 8'sb11111111, 8'sb00001010, 8'sb00010001, 8'sb00100001, 8'sb00001111, 8'sb00010000, 8'sb00001011, 8'sb11111111, 8'sb11111010, 8'sb00001000, 8'sb00001110, 8'sb11111111, 8'sb00001111, 8'sb00010001, 8'sb00000000, 8'sb00000001, 8'sb00000111, 8'sb00010100, 8'sb00001110, 8'sb00001111, 8'sb00001101, 8'sb00001011, 8'sb00011010, 8'sb00010100, 8'sb00111001, 8'sb00011100, 8'sb11111110, 8'sb11111100, 8'sb00000010, 8'sb00000111, 8'sb00011001, 8'sb00001111, 8'sb00001100, 8'sb00010000, 8'sb00001110, 8'sb00011110, 8'sb00100001, 8'sb00110000, 8'sb00101011, 8'sb00001111, 8'sb00000110, 8'sb00011000, 8'sb00010101, 8'sb00010100, 8'sb00100110, 8'sb00010110, 8'sb00001100, 8'sb00010000, 8'sb00010010, 8'sb00011000, 8'sb00100011, 8'sb00010100, 8'sb00000110, 8'sb00001110, 8'sb00011010, 8'sb00011100, 8'sb00011010, 8'sb00011110, 8'sb00011111, 8'sb00010001, 8'sb00001100, 8'sb00010000, 8'sb00001110, 8'sb00011111, 8'sb00100010, 8'sb00000011, 8'sb00000001, 8'sb00010010, 8'sb00011101, 8'sb00011000, 8'sb00001110, 8'sb00010010, 8'sb00010100, 8'sb00001011, 8'sb00001011, 8'sb00010000, 8'sb00010000, 8'sb00010111, 8'sb00010110, 8'sb00010111, 8'sb00011010, 8'sb00011101, 8'sb00011101, 8'sb00010111, 8'sb00010011, 8'sb00001101, 8'sb00001111, 8'sb00001100, 8'sb00010000, 8'sb00001101, 8'sb00001100, 8'sb00001100, 8'sb00001011, 8'sb00001001, 8'sb00001101, 8'sb00001101, 8'sb00001000, 8'sb00001110, 8'sb00010110, 8'sb00001110, 8'sb00000011, 8'sb00001110, 8'sb00001101, 8'sb00001111, 8'sb00001101, 8'sb00001100, 8'sb11111111, 8'sb11110010, 8'sb11111010, 8'sb11111110, 8'sb00001000, 8'sb00001000, 8'sb00000110, 8'sb00000100, 8'sb00001001, 8'sb00001101, 8'sb00001111, 8'sb00001111, 8'sb00001100, 8'sb00001110, 8'sb00000111, 8'sb00000111, 8'sb00000010, 8'sb11111111, 8'sb11111010, 8'sb11111111, 8'sb00000001, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00001100,
    8'sb00001111, 8'sb00001100, 8'sb00001111, 8'sb00010000, 8'sb00001100, 8'sb00001110, 8'sb00001101, 8'sb00010001, 8'sb00001110, 8'sb00010000, 8'sb00001101, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00001110, 8'sb00001010, 8'sb00001000, 8'sb00001001, 8'sb00001010, 8'sb00000111, 8'sb00001100, 8'sb00010000, 8'sb00010000, 8'sb00010000, 8'sb00010000, 8'sb00001101, 8'sb00001101, 8'sb00001101, 8'sb00001111, 8'sb00010010, 8'sb00001110, 8'sb00010010, 8'sb00010100, 8'sb00001110, 8'sb00000110, 8'sb00010000, 8'sb00001111, 8'sb00001110, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00010110, 8'sb00011000, 8'sb00010001, 8'sb00000011, 8'sb00011010, 8'sb00100010, 8'sb00010001, 8'sb00000101, 8'sb00001100, 8'sb00010001, 8'sb00001111, 8'sb00001100, 8'sb00010100, 8'sb00011111, 8'sb00011001, 8'sb00011000, 8'sb00001110, 8'sb00001000, 8'sb00100100, 8'sb00011100, 8'sb00010010, 8'sb00001101, 8'sb00000100, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00011001, 8'sb00011011, 8'sb00001111, 8'sb00001101, 8'sb11101010, 8'sb00011011, 8'sb00100100, 8'sb00001011, 8'sb00001100, 8'sb00001111, 8'sb00001001, 8'sb00010000, 8'sb00001110, 8'sb00001101, 8'sb00010010, 8'sb11111011, 8'sb11110011, 8'sb11100110, 8'sb11111110, 8'sb00110010, 8'sb00010011, 8'sb00011100, 8'sb00101011, 8'sb00001111, 8'sb00010001, 8'sb00010000, 8'sb00001101, 8'sb00001101, 8'sb00000100, 8'sb11110011, 8'sb11111001, 8'sb00010000, 8'sb00100111, 8'sb00100100, 8'sb00011100, 8'sb00011111, 8'sb00001011, 8'sb11110110, 8'sb00001010, 8'sb00001110, 8'sb00010001, 8'sb00001011, 8'sb00000101, 8'sb00001011, 8'sb00011100, 8'sb00010111, 8'sb00100100, 8'sb00100000, 8'sb00011001, 8'sb00000110, 8'sb00000000, 8'sb11111011, 8'sb00001110, 8'sb00001101, 8'sb00001111, 8'sb00001100, 8'sb11111101, 8'sb00000000, 8'sb00001000, 8'sb00000000, 8'sb00010001, 8'sb00001100, 8'sb00000000, 8'sb00000110, 8'sb00001001, 8'sb00001010, 8'sb00010010, 8'sb00001101, 8'sb00001101, 8'sb00001111, 8'sb00010011, 8'sb00001111, 8'sb00001011, 8'sb00000001, 8'sb00000001, 8'sb00001000, 8'sb00000110, 8'sb00000101, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00001100, 8'sb00010001, 8'sb00010000, 8'sb00010111, 8'sb00011000, 8'sb00001110, 8'sb00001000, 8'sb00001011, 8'sb00001101, 8'sb00000111, 8'sb00001001, 8'sb00010110, 8'sb00010101, 8'sb00010010, 8'sb00001100, 8'sb00001110, 8'sb00001111, 8'sb00010001, 8'sb00010100, 8'sb00001110, 8'sb00000110, 8'sb00001100, 8'sb00001110, 8'sb00001100, 8'sb00010001, 8'sb00010111, 8'sb00010010, 8'sb00010001, 8'sb00001110, 8'sb00001110, 8'sb00001111, 8'sb00010010, 8'sb00001111, 8'sb00010011, 8'sb00010010, 8'sb00010100, 8'sb00010111, 8'sb00001111, 8'sb00001110, 8'sb00001111, 8'sb00010000, 8'sb00010001, 8'sb00001100,
    8'sb00010000, 8'sb00001101, 8'sb00001110, 8'sb00001101, 8'sb00001111, 8'sb00001100, 8'sb00001101, 8'sb00001101, 8'sb00010000, 8'sb00001111, 8'sb00001100, 8'sb00001111, 8'sb00010000, 8'sb00001011, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00010111, 8'sb00011100, 8'sb00100010, 8'sb00100010, 8'sb00011010, 8'sb00011000, 8'sb00010011, 8'sb00010100, 8'sb00001111, 8'sb00010000, 8'sb00001110, 8'sb00001111, 8'sb00010001, 8'sb00010011, 8'sb00010001, 8'sb00001010, 8'sb00010100, 8'sb00010111, 8'sb00001010, 8'sb00000101, 8'sb00010011, 8'sb00001111, 8'sb00010000, 8'sb00001100, 8'sb00001111, 8'sb00001110, 8'sb00001111, 8'sb00000000, 8'sb00000111, 8'sb00000000, 8'sb00001001, 8'sb00101000, 8'sb00011110, 8'sb11111000, 8'sb00000100, 8'sb11111000, 8'sb00000111, 8'sb00001101, 8'sb00001011, 8'sb00001100, 8'sb00001111, 8'sb00010001, 8'sb00001101, 8'sb11111111, 8'sb00000010, 8'sb00110001, 8'sb00000011, 8'sb11111011, 8'sb00001111, 8'sb11110010, 8'sb11110100, 8'sb00001110, 8'sb00001100, 8'sb00010001, 8'sb00010010, 8'sb00010010, 8'sb11111110, 8'sb11111000, 8'sb11101111, 8'sb01000001, 8'sb00000111, 8'sb00001011, 8'sb00001001, 8'sb00001010, 8'sb00000110, 8'sb00001110, 8'sb00001100, 8'sb00010000, 8'sb00010100, 8'sb00000101, 8'sb00010011, 8'sb00000110, 8'sb11110010, 8'sb00111000, 8'sb00010100, 8'sb00010101, 8'sb00001010, 8'sb00011110, 8'sb00010101, 8'sb00001111, 8'sb00001100, 8'sb00010010, 8'sb00000101, 8'sb00010001, 8'sb00001100, 8'sb00000111, 8'sb00001111, 8'sb00100111, 8'sb00010101, 8'sb00010000, 8'sb00010110, 8'sb00001101, 8'sb00010010, 8'sb00001100, 8'sb00001111, 8'sb00010011, 8'sb00001011, 8'sb00011010, 8'sb00010001, 8'sb00010000, 8'sb00010110, 8'sb00011110, 8'sb00010001, 8'sb00010000, 8'sb00001110, 8'sb00000110, 8'sb00001100, 8'sb00001101, 8'sb00001101, 8'sb00010010, 8'sb00001010, 8'sb00000100, 8'sb00001011, 8'sb00001100, 8'sb00010100, 8'sb00010111, 8'sb00010110, 8'sb00010101, 8'sb00001110, 8'sb00001010, 8'sb00001010, 8'sb00001101, 8'sb00001100, 8'sb00010010, 8'sb00010010, 8'sb00010011, 8'sb00000101, 8'sb00000011, 8'sb00010111, 8'sb00011111, 8'sb00010110, 8'sb00010000, 8'sb00000001, 8'sb11111110, 8'sb00001100, 8'sb00001110, 8'sb00001101, 8'sb00010000, 8'sb00010001, 8'sb00000110, 8'sb11111111, 8'sb11111111, 8'sb00000010, 8'sb00010010, 8'sb00001111, 8'sb00001001, 8'sb00001010, 8'sb00001100, 8'sb00001111, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00010000, 8'sb00010111, 8'sb00010100, 8'sb00011001, 8'sb00001001, 8'sb00001100, 8'sb00010100, 8'sb00011101, 8'sb00100001, 8'sb00010010, 8'sb00001101, 8'sb00001110, 8'sb00001101, 8'sb00001111, 8'sb00001111, 8'sb00010001, 8'sb00011000, 8'sb00011000, 8'sb00010111, 8'sb00011000, 8'sb00010100, 8'sb00010000, 8'sb00010000, 8'sb00010000, 8'sb00001101, 8'sb00001111,
    8'sb00010011, 8'sb00010001, 8'sb00010011, 8'sb00010011, 8'sb00010001, 8'sb00010010, 8'sb00010100, 8'sb00010101, 8'sb00010011, 8'sb00010010, 8'sb00010001, 8'sb00010001, 8'sb00010011, 8'sb00010010, 8'sb00010000, 8'sb00010010, 8'sb00010000, 8'sb00010100, 8'sb00010011, 8'sb00010110, 8'sb00011000, 8'sb00011001, 8'sb00010100, 8'sb00010111, 8'sb00010110, 8'sb00010101, 8'sb00010010, 8'sb00010100, 8'sb00010100, 8'sb00010010, 8'sb00010001, 8'sb00001110, 8'sb00000100, 8'sb11111111, 8'sb00000001, 8'sb00000010, 8'sb00000101, 8'sb00011011, 8'sb00010110, 8'sb00011101, 8'sb00010001, 8'sb00010000, 8'sb00010010, 8'sb00001110, 8'sb00001011, 8'sb11111010, 8'sb11110001, 8'sb00000110, 8'sb00001011, 8'sb00010001, 8'sb00000101, 8'sb00010001, 8'sb00000100, 8'sb00001000, 8'sb00001110, 8'sb00010000, 8'sb00010011, 8'sb00001111, 8'sb11111010, 8'sb11101100, 8'sb00000101, 8'sb00001110, 8'sb00001110, 8'sb00001001, 8'sb00001010, 8'sb11111011, 8'sb11110100, 8'sb00000000, 8'sb00001010, 8'sb00010001, 8'sb00010000, 8'sb00001011, 8'sb11111001, 8'sb00001100, 8'sb00011101, 8'sb00011111, 8'sb00011010, 8'sb00001110, 8'sb11110110, 8'sb00000000, 8'sb00001000, 8'sb00010100, 8'sb00001000, 8'sb00010000, 8'sb00010000, 8'sb00001100, 8'sb00010001, 8'sb00101000, 8'sb00011110, 8'sb00001110, 8'sb00010011, 8'sb00011010, 8'sb00010010, 8'sb00010100, 8'sb00010101, 8'sb00101100, 8'sb00011010, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00001110, 8'sb00100011, 8'sb00011001, 8'sb00001100, 8'sb00001000, 8'sb00011110, 8'sb00011000, 8'sb11111111, 8'sb00001110, 8'sb00010011, 8'sb00001110, 8'sb00001101, 8'sb00010100, 8'sb00001101, 8'sb11111011, 8'sb00001010, 8'sb00011100, 8'sb00100010, 8'sb00010011, 8'sb00011111, 8'sb00000010, 8'sb00000101, 8'sb00000001, 8'sb00000110, 8'sb00001000, 8'sb00010001, 8'sb00010011, 8'sb00001101, 8'sb11111101, 8'sb11111000, 8'sb11111110, 8'sb00001101, 8'sb00011000, 8'sb00001111, 8'sb00000101, 8'sb00000101, 8'sb00001111, 8'sb00001100, 8'sb00000100, 8'sb00010010, 8'sb00001111, 8'sb00010001, 8'sb00000100, 8'sb00001000, 8'sb00001110, 8'sb00011000, 8'sb00011001, 8'sb00011010, 8'sb00010100, 8'sb00001010, 8'sb00001101, 8'sb00001001, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00010000, 8'sb00001110, 8'sb00000100, 8'sb00011010, 8'sb00001111, 8'sb00010001, 8'sb00001101, 8'sb00010111, 8'sb00000110, 8'sb00000111, 8'sb00001101, 8'sb00010001, 8'sb00010000, 8'sb00010010, 8'sb00010100, 8'sb00010101, 8'sb00010000, 8'sb00010001, 8'sb00001010, 8'sb00000100, 8'sb00000101, 8'sb00001101, 8'sb00001110, 8'sb00010101, 8'sb00010110, 8'sb00010010, 8'sb00010001, 8'sb00010011, 8'sb00010100, 8'sb00010001, 8'sb00010101, 8'sb00010011, 8'sb00010100, 8'sb00010101, 8'sb00010101, 8'sb00010001, 8'sb00001111, 8'sb00010001, 8'sb00010011, 8'sb00010001, 8'sb00010100,
    8'sb00001010, 8'sb00001101, 8'sb00001011, 8'sb00001001, 8'sb00001011, 8'sb00001010, 8'sb00001011, 8'sb00001011, 8'sb00001000, 8'sb00001011, 8'sb00001100, 8'sb00001010, 8'sb00001011, 8'sb00001100, 8'sb00001001, 8'sb00001101, 8'sb00001000, 8'sb00001010, 8'sb00001100, 8'sb00001010, 8'sb11111111, 8'sb00000000, 8'sb00001011, 8'sb00010001, 8'sb00001110, 8'sb00001011, 8'sb00001001, 8'sb00001011, 8'sb00001001, 8'sb00001001, 8'sb00001000, 8'sb00000101, 8'sb00001010, 8'sb00001000, 8'sb00001100, 8'sb00001011, 8'sb00010101, 8'sb00011011, 8'sb00011001, 8'sb00010110, 8'sb00001110, 8'sb00001011, 8'sb00001010, 8'sb00001010, 8'sb00000100, 8'sb00010000, 8'sb00010000, 8'sb00001101, 8'sb00010000, 8'sb00001110, 8'sb00010111, 8'sb00010011, 8'sb00101111, 8'sb00101111, 8'sb00010100, 8'sb00001110, 8'sb00001010, 8'sb00001000, 8'sb00000001, 8'sb00001001, 8'sb00011000, 8'sb00011101, 8'sb00010010, 8'sb11110011, 8'sb11110010, 8'sb00010000, 8'sb00111111, 8'sb00110100, 8'sb00011001, 8'sb00001011, 8'sb00001001, 8'sb00001000, 8'sb00010000, 8'sb00100000, 8'sb00100100, 8'sb00000101, 8'sb00000100, 8'sb11101001, 8'sb00001011, 8'sb00101100, 8'sb00110011, 8'sb00011100, 8'sb00010010, 8'sb00001010, 8'sb00001101, 8'sb00001100, 8'sb00011000, 8'sb00011010, 8'sb00001000, 8'sb00010001, 8'sb11111101, 8'sb00000011, 8'sb00011101, 8'sb00101001, 8'sb00100000, 8'sb00010000, 8'sb00001010, 8'sb00001011, 8'sb00001000, 8'sb00001101, 8'sb00010000, 8'sb00010000, 8'sb00001001, 8'sb00010100, 8'sb00001010, 8'sb00001111, 8'sb00011100, 8'sb00011000, 8'sb00001000, 8'sb00001100, 8'sb00010000, 8'sb00001011, 8'sb00001000, 8'sb00001010, 8'sb00010010, 8'sb00010010, 8'sb00001001, 8'sb00001001, 8'sb00010011, 8'sb00011001, 8'sb00011101, 8'sb00001101, 8'sb00001000, 8'sb11111111, 8'sb00001111, 8'sb00001001, 8'sb00001010, 8'sb00000111, 8'sb00010011, 8'sb00010010, 8'sb00010011, 8'sb00010011, 8'sb00001011, 8'sb00001111, 8'sb00000101, 8'sb00001000, 8'sb00000100, 8'sb00000100, 8'sb00001110, 8'sb00001100, 8'sb00001001, 8'sb00001001, 8'sb00010100, 8'sb00010111, 8'sb00010100, 8'sb00010100, 8'sb00011010, 8'sb00001110, 8'sb00001100, 8'sb00001111, 8'sb00010101, 8'sb00011011, 8'sb00001101, 8'sb00001011, 8'sb00001011, 8'sb00000110, 8'sb00001000, 8'sb00010011, 8'sb00001100, 8'sb00001010, 8'sb00010010, 8'sb00011000, 8'sb00001001, 8'sb00000001, 8'sb00010110, 8'sb00010000, 8'sb00001101, 8'sb00001010, 8'sb00001001, 8'sb00001001, 8'sb00000101, 8'sb00000100, 8'sb00000101, 8'sb00001111, 8'sb00001111, 8'sb00010000, 8'sb00001110, 8'sb00010010, 8'sb00010000, 8'sb00001010, 8'sb00001000, 8'sb00001011, 8'sb00001000, 8'sb00001100, 8'sb00001000, 8'sb00001010, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00001110, 8'sb00001011, 8'sb00001010, 8'sb00001010, 8'sb00001101, 8'sb00001010, 8'sb00001010,
    8'sb00001110, 8'sb00001111, 8'sb00001111, 8'sb00001011, 8'sb00001011, 8'sb00001110, 8'sb00001111, 8'sb00001111, 8'sb00001111, 8'sb00001011, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00001100, 8'sb00001110, 8'sb00001011, 8'sb00001101, 8'sb00010011, 8'sb00010100, 8'sb00010111, 8'sb00011011, 8'sb00011000, 8'sb00001100, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00001001, 8'sb00000110, 8'sb00001110, 8'sb00010000, 8'sb00010100, 8'sb00011011, 8'sb00010100, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00010010, 8'sb00001110, 8'sb00001100, 8'sb00001100, 8'sb00001011, 8'sb11111101, 8'sb00001001, 8'sb00001111, 8'sb00000111, 8'sb00000011, 8'sb00010111, 8'sb00011101, 8'sb00000101, 8'sb00001001, 8'sb00001110, 8'sb00011100, 8'sb00001100, 8'sb00001111, 8'sb00001010, 8'sb11111100, 8'sb11111110, 8'sb00000000, 8'sb00001011, 8'sb00001111, 8'sb00010101, 8'sb00000100, 8'sb00000110, 8'sb00001001, 8'sb00100100, 8'sb00101111, 8'sb00001100, 8'sb00001011, 8'sb00001011, 8'sb00010000, 8'sb00100000, 8'sb00101000, 8'sb00101001, 8'sb00110010, 8'sb00001101, 8'sb11110000, 8'sb00000011, 8'sb00010111, 8'sb00100110, 8'sb00011100, 8'sb00001111, 8'sb00001100, 8'sb00001101, 8'sb00011100, 8'sb00101110, 8'sb00100100, 8'sb00011010, 8'sb00011110, 8'sb00011010, 8'sb00001000, 8'sb00001001, 8'sb00010100, 8'sb00011001, 8'sb00001110, 8'sb00001110, 8'sb00001100, 8'sb00001010, 8'sb00001010, 8'sb00000111, 8'sb00010001, 8'sb00001110, 8'sb00010110, 8'sb11111111, 8'sb00000111, 8'sb00000001, 8'sb00000001, 8'sb00010110, 8'sb00001100, 8'sb00001100, 8'sb00001100, 8'sb00000110, 8'sb00000110, 8'sb00001011, 8'sb00010110, 8'sb00011010, 8'sb00001000, 8'sb11111101, 8'sb00000011, 8'sb11111111, 8'sb00000101, 8'sb00010000, 8'sb00001110, 8'sb00001110, 8'sb00001011, 8'sb00001001, 8'sb00000111, 8'sb00001101, 8'sb00010011, 8'sb00100111, 8'sb00010011, 8'sb11111110, 8'sb00010011, 8'sb00010100, 8'sb00010100, 8'sb00010110, 8'sb00001010, 8'sb00001110, 8'sb00001101, 8'sb00001000, 8'sb00000110, 8'sb00000110, 8'sb00001110, 8'sb00010111, 8'sb00011010, 8'sb00000010, 8'sb00000111, 8'sb00000111, 8'sb00001100, 8'sb00010111, 8'sb00001101, 8'sb00001011, 8'sb00001011, 8'sb00001010, 8'sb00000111, 8'sb00000101, 8'sb00010001, 8'sb00011011, 8'sb00100010, 8'sb00001011, 8'sb00000110, 8'sb00000000, 8'sb00001011, 8'sb00001101, 8'sb00001001, 8'sb00001101, 8'sb00001010, 8'sb00001101, 8'sb00000111, 8'sb00001001, 8'sb00010100, 8'sb00011001, 8'sb00011101, 8'sb00010010, 8'sb00010110, 8'sb00010010, 8'sb00001101, 8'sb00001010, 8'sb00001011, 8'sb00001111, 8'sb00001011, 8'sb00001110, 8'sb00001100, 8'sb00001011, 8'sb00001101, 8'sb00010001, 8'sb00010101, 8'sb00010001, 8'sb00001111, 8'sb00001101, 8'sb00001101, 8'sb00001101, 8'sb00001100, 8'sb00001110,
    8'sb00010011, 8'sb00010011, 8'sb00010011, 8'sb00001110, 8'sb00010000, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00010001, 8'sb00010001, 8'sb00010001, 8'sb00010000, 8'sb00010000, 8'sb00010010, 8'sb00010011, 8'sb00010000, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00010001, 8'sb00010011, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00001101, 8'sb00001101, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00010001, 8'sb00010001, 8'sb00001111, 8'sb00001010, 8'sb00001100, 8'sb00010011, 8'sb00011000, 8'sb00100100, 8'sb00010110, 8'sb00010010, 8'sb00000100, 8'sb00010011, 8'sb00010100, 8'sb00010000, 8'sb00010010, 8'sb00010001, 8'sb00001001, 8'sb00000100, 8'sb00001110, 8'sb00000110, 8'sb00001100, 8'sb00011110, 8'sb00011101, 8'sb00010110, 8'sb00001110, 8'sb00000111, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00010001, 8'sb00010100, 8'sb00010110, 8'sb00001111, 8'sb00010010, 8'sb11111111, 8'sb00001010, 8'sb00110101, 8'sb00011000, 8'sb00011010, 8'sb11110011, 8'sb00001100, 8'sb00010000, 8'sb00001011, 8'sb00001110, 8'sb00001111, 8'sb00010111, 8'sb00001010, 8'sb00000111, 8'sb11011000, 8'sb00101010, 8'sb00101111, 8'sb00011110, 8'sb00011111, 8'sb11110011, 8'sb00001010, 8'sb00001111, 8'sb00001111, 8'sb00001000, 8'sb00001011, 8'sb00001000, 8'sb11111110, 8'sb00000001, 8'sb00000111, 8'sb00100110, 8'sb00100100, 8'sb00100111, 8'sb01000001, 8'sb00110010, 8'sb00001110, 8'sb00010010, 8'sb00001110, 8'sb00010101, 8'sb00011101, 8'sb00000010, 8'sb00001000, 8'sb00001111, 8'sb00010101, 8'sb00010100, 8'sb00010010, 8'sb00001001, 8'sb00001111, 8'sb00011010, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00010110, 8'sb00011101, 8'sb00001010, 8'sb00010111, 8'sb00001101, 8'sb00011000, 8'sb00001000, 8'sb00001011, 8'sb00001010, 8'sb00001011, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00000100, 8'sb00000100, 8'sb00010100, 8'sb00010100, 8'sb00001100, 8'sb00001001, 8'sb00001000, 8'sb00000111, 8'sb00000000, 8'sb11111110, 8'sb00001110, 8'sb00010010, 8'sb00001111, 8'sb00010010, 8'sb00001101, 8'sb00011100, 8'sb00001101, 8'sb00010001, 8'sb00010010, 8'sb00010011, 8'sb00000100, 8'sb00000110, 8'sb00000010, 8'sb11111111, 8'sb00001110, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00001000, 8'sb00010101, 8'sb00001000, 8'sb00001100, 8'sb00010110, 8'sb00001110, 8'sb00000100, 8'sb00001011, 8'sb00001011, 8'sb00001110, 8'sb00010100, 8'sb00010000, 8'sb00010010, 8'sb00001111, 8'sb00001101, 8'sb00001011, 8'sb00001001, 8'sb00010001, 8'sb00010001, 8'sb00010011, 8'sb00010000, 8'sb00010001, 8'sb00001100, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00010001, 8'sb00010001, 8'sb00001110, 8'sb00010010, 8'sb00010001, 8'sb00010000, 8'sb00001110, 8'sb00001011, 8'sb00001110, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00010000,
    8'sb00010001, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00001100, 8'sb00001011, 8'sb00001010, 8'sb00001011, 8'sb00001011, 8'sb00001001, 8'sb00001110, 8'sb00010010, 8'sb00010001, 8'sb00001101, 8'sb00001101, 8'sb00010000, 8'sb00001101, 8'sb00001010, 8'sb00000000, 8'sb00000010, 8'sb00001001, 8'sb00001001, 8'sb00000110, 8'sb00001111, 8'sb00010000, 8'sb00010111, 8'sb00100010, 8'sb00010010, 8'sb00010001, 8'sb00001110, 8'sb00001101, 8'sb00000001, 8'sb00000110, 8'sb00010100, 8'sb00011011, 8'sb00011010, 8'sb00001000, 8'sb00001001, 8'sb00010000, 8'sb00001101, 8'sb00011001, 8'sb00011000, 8'sb00001110, 8'sb00010000, 8'sb00001100, 8'sb00000000, 8'sb00001011, 8'sb00010001, 8'sb00100000, 8'sb00001100, 8'sb00001110, 8'sb00010110, 8'sb00010101, 8'sb00010001, 8'sb00001110, 8'sb00011011, 8'sb00001111, 8'sb00010000, 8'sb00001101, 8'sb00010001, 8'sb00011000, 8'sb00010111, 8'sb00101110, 8'sb00001001, 8'sb11110001, 8'sb00010110, 8'sb00000100, 8'sb00000100, 8'sb00000101, 8'sb00001110, 8'sb00001111, 8'sb00001111, 8'sb00010001, 8'sb00011110, 8'sb00101100, 8'sb00100000, 8'sb00100001, 8'sb11111111, 8'sb11110100, 8'sb00010110, 8'sb00011100, 8'sb00010110, 8'sb00010110, 8'sb00001011, 8'sb00001101, 8'sb00010001, 8'sb00010000, 8'sb00100000, 8'sb00100011, 8'sb00010111, 8'sb00010001, 8'sb11111111, 8'sb11101000, 8'sb00010111, 8'sb00001101, 8'sb00010001, 8'sb00010111, 8'sb00010010, 8'sb00001101, 8'sb00001101, 8'sb00001010, 8'sb00010111, 8'sb00010110, 8'sb00001101, 8'sb00001100, 8'sb11110000, 8'sb11111101, 8'sb00011100, 8'sb00010010, 8'sb00010100, 8'sb00000010, 8'sb00001100, 8'sb00001101, 8'sb00001111, 8'sb00000111, 8'sb00001111, 8'sb00001111, 8'sb00001001, 8'sb00000000, 8'sb11101100, 8'sb00010101, 8'sb00001110, 8'sb00001110, 8'sb00000110, 8'sb11111110, 8'sb00001010, 8'sb00001100, 8'sb00010001, 8'sb00001100, 8'sb00010110, 8'sb00001111, 8'sb11111111, 8'sb11111100, 8'sb00010100, 8'sb00010011, 8'sb00001110, 8'sb00001010, 8'sb00000010, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010001, 8'sb00001011, 8'sb00001001, 8'sb00000100, 8'sb00000100, 8'sb00000101, 8'sb00011001, 8'sb00010011, 8'sb00010011, 8'sb00010001, 8'sb00010100, 8'sb00010100, 8'sb00001111, 8'sb00001101, 8'sb00010001, 8'sb00001100, 8'sb00001110, 8'sb00001000, 8'sb00001011, 8'sb00001101, 8'sb00001111, 8'sb00010001, 8'sb00010100, 8'sb00010100, 8'sb00010111, 8'sb00010001, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00001101, 8'sb00010001, 8'sb00010001, 8'sb00010010, 8'sb00010101, 8'sb00010011, 8'sb00010011, 8'sb00010011, 8'sb00010011, 8'sb00001110, 8'sb00010010, 8'sb00010000, 8'sb00010001,
    8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00001011, 8'sb00001010, 8'sb00001010, 8'sb00001100, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00001110, 8'sb00001011, 8'sb00001010, 8'sb00001110, 8'sb00001100, 8'sb00001110, 8'sb00001100, 8'sb00001111, 8'sb00001101, 8'sb00001100, 8'sb00010010, 8'sb00001111, 8'sb00001100, 8'sb00000110, 8'sb00001000, 8'sb00001100, 8'sb00001010, 8'sb00001010, 8'sb00001101, 8'sb00001110, 8'sb00001101, 8'sb00001110, 8'sb00010010, 8'sb00010001, 8'sb00001001, 8'sb00000111, 8'sb11110111, 8'sb00001100, 8'sb11111111, 8'sb11111101, 8'sb00001100, 8'sb00001100, 8'sb00001011, 8'sb00001101, 8'sb00001010, 8'sb00001001, 8'sb00010010, 8'sb00011000, 8'sb00101101, 8'sb00100100, 8'sb00100101, 8'sb00100101, 8'sb00100101, 8'sb11111101, 8'sb00000011, 8'sb00001010, 8'sb00001101, 8'sb00001010, 8'sb00000001, 8'sb00001001, 8'sb00010101, 8'sb00010100, 8'sb00100011, 8'sb00110111, 8'sb00101010, 8'sb00011000, 8'sb00010000, 8'sb00011011, 8'sb00001110, 8'sb00001011, 8'sb00001101, 8'sb00001111, 8'sb00001100, 8'sb00011010, 8'sb00010111, 8'sb00011110, 8'sb00101001, 8'sb00011110, 8'sb00010110, 8'sb00011001, 8'sb00011011, 8'sb00100011, 8'sb00011000, 8'sb00001011, 8'sb00001100, 8'sb00010011, 8'sb00011111, 8'sb00010100, 8'sb00010101, 8'sb00000110, 8'sb11101010, 8'sb00000110, 8'sb00001110, 8'sb00010010, 8'sb00010000, 8'sb00001111, 8'sb00000101, 8'sb00001101, 8'sb00001110, 8'sb00001110, 8'sb00010001, 8'sb00001011, 8'sb00000010, 8'sb00000001, 8'sb11110101, 8'sb11110111, 8'sb00000100, 8'sb11111101, 8'sb00001101, 8'sb11111101, 8'sb00000100, 8'sb00001100, 8'sb00001100, 8'sb00001101, 8'sb00001100, 8'sb11111101, 8'sb00000011, 8'sb00011000, 8'sb11111100, 8'sb11101110, 8'sb00000001, 8'sb00000110, 8'sb11111010, 8'sb11111100, 8'sb00000101, 8'sb00001010, 8'sb00001110, 8'sb00000111, 8'sb00001100, 8'sb00001100, 8'sb00010010, 8'sb00001100, 8'sb11111100, 8'sb00001001, 8'sb00001001, 8'sb00011001, 8'sb00010110, 8'sb00001111, 8'sb00000111, 8'sb00001101, 8'sb00001010, 8'sb00001011, 8'sb00010011, 8'sb00010101, 8'sb00010100, 8'sb11111010, 8'sb00000010, 8'sb00001001, 8'sb00001000, 8'sb00010001, 8'sb00010101, 8'sb00010110, 8'sb00001110, 8'sb00001010, 8'sb00001101, 8'sb00001011, 8'sb00001111, 8'sb00011010, 8'sb00011110, 8'sb00001100, 8'sb00001000, 8'sb00000000, 8'sb11111100, 8'sb11110111, 8'sb00000011, 8'sb00011010, 8'sb00001110, 8'sb00001011, 8'sb00001011, 8'sb00001011, 8'sb00010001, 8'sb00011110, 8'sb00100010, 8'sb00011101, 8'sb00011111, 8'sb00100010, 8'sb00100110, 8'sb00100010, 8'sb00010101, 8'sb00010110, 8'sb00001111, 8'sb00001011, 8'sb00001101, 8'sb00001110, 8'sb00001111, 8'sb00010100, 8'sb00011000, 8'sb00011011, 8'sb00100000, 8'sb00100100, 8'sb00100001, 8'sb00011010, 8'sb00010000, 8'sb00001111, 8'sb00001100, 8'sb00001100,
    8'sb00010100, 8'sb00010000, 8'sb00001111, 8'sb00010011, 8'sb00010011, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00010010, 8'sb00010000, 8'sb00010000, 8'sb00010001, 8'sb00010011, 8'sb00010001, 8'sb00010100, 8'sb00010100, 8'sb00010010, 8'sb00010000, 8'sb00001111, 8'sb00001100, 8'sb00001001, 8'sb00001001, 8'sb00001110, 8'sb00010101, 8'sb00010100, 8'sb00010111, 8'sb00010001, 8'sb00010001, 8'sb00010010, 8'sb00010010, 8'sb00010100, 8'sb00010011, 8'sb00001010, 8'sb00000010, 8'sb00000110, 8'sb00010000, 8'sb00000111, 8'sb00001101, 8'sb00011010, 8'sb00011011, 8'sb00001110, 8'sb00010010, 8'sb00010011, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00000100, 8'sb11111111, 8'sb11110010, 8'sb11100111, 8'sb11101011, 8'sb00000010, 8'sb00001101, 8'sb00010100, 8'sb00001100, 8'sb00001110, 8'sb00001111, 8'sb00010000, 8'sb00010001, 8'sb00000011, 8'sb11111000, 8'sb11101101, 8'sb11110101, 8'sb00000000, 8'sb00010010, 8'sb00000100, 8'sb00000110, 8'sb11111000, 8'sb11111000, 8'sb00001011, 8'sb00010011, 8'sb00010010, 8'sb00001110, 8'sb00010001, 8'sb00100001, 8'sb00110110, 8'sb00111111, 8'sb00011010, 8'sb00000101, 8'sb00000110, 8'sb00010011, 8'sb00000010, 8'sb11111101, 8'sb00001111, 8'sb00010000, 8'sb00010000, 8'sb00011011, 8'sb00100111, 8'sb00101010, 8'sb00011010, 8'sb00001011, 8'sb00010001, 8'sb00010011, 8'sb00001101, 8'sb00001111, 8'sb00011011, 8'sb00010011, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00011100, 8'sb00010110, 8'sb00001100, 8'sb00000111, 8'sb00011001, 8'sb00010110, 8'sb00001111, 8'sb00010010, 8'sb00010110, 8'sb00011010, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00001100, 8'sb11111011, 8'sb00001110, 8'sb00011011, 8'sb00010111, 8'sb00011010, 8'sb00010001, 8'sb00001000, 8'sb00010010, 8'sb00010011, 8'sb00000100, 8'sb11111111, 8'sb00001111, 8'sb00010010, 8'sb00001101, 8'sb11110011, 8'sb11101010, 8'sb00010010, 8'sb00010111, 8'sb00011100, 8'sb00001111, 8'sb00001100, 8'sb00010010, 8'sb00001100, 8'sb00000000, 8'sb00000000, 8'sb00010001, 8'sb00010010, 8'sb00001100, 8'sb00000000, 8'sb11111101, 8'sb00000001, 8'sb00001010, 8'sb00010011, 8'sb00011000, 8'sb00010110, 8'sb00010100, 8'sb00000010, 8'sb11111111, 8'sb00001101, 8'sb00010011, 8'sb00001111, 8'sb00010001, 8'sb00010100, 8'sb00010100, 8'sb00001111, 8'sb00001111, 8'sb00010100, 8'sb00011001, 8'sb00010111, 8'sb00011000, 8'sb00001000, 8'sb00000110, 8'sb00001101, 8'sb00010001, 8'sb00010010, 8'sb00010000, 8'sb00010010, 8'sb00001111, 8'sb00001100, 8'sb00010100, 8'sb00001010, 8'sb00001001, 8'sb00000110, 8'sb00001001, 8'sb00001001, 8'sb00001110, 8'sb00001101, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00010000, 8'sb00001111, 8'sb00001010, 8'sb00000101, 8'sb00001000, 8'sb00001100, 8'sb00001100, 8'sb00010001, 8'sb00010010, 8'sb00001111,
    8'sb00010011, 8'sb00010000, 8'sb00010000, 8'sb00010001, 8'sb00010000, 8'sb00010010, 8'sb00010000, 8'sb00010011, 8'sb00001111, 8'sb00010001, 8'sb00010010, 8'sb00010010, 8'sb00010011, 8'sb00010001, 8'sb00010010, 8'sb00001111, 8'sb00010001, 8'sb00010010, 8'sb00010001, 8'sb00010010, 8'sb00010101, 8'sb00010110, 8'sb00011010, 8'sb00010011, 8'sb00010010, 8'sb00010100, 8'sb00010001, 8'sb00010010, 8'sb00010100, 8'sb00010011, 8'sb00010100, 8'sb00001110, 8'sb00001111, 8'sb00001011, 8'sb00001001, 8'sb00001000, 8'sb11111110, 8'sb00000101, 8'sb00010000, 8'sb00010011, 8'sb00001010, 8'sb00010011, 8'sb00010000, 8'sb00001110, 8'sb00001001, 8'sb11111001, 8'sb11110101, 8'sb11111110, 8'sb11111100, 8'sb00001010, 8'sb00000101, 8'sb00000100, 8'sb00001001, 8'sb00000110, 8'sb00000110, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb11111010, 8'sb11110110, 8'sb11110101, 8'sb00000010, 8'sb00010000, 8'sb00010001, 8'sb11111011, 8'sb00000101, 8'sb00001000, 8'sb11111001, 8'sb11111110, 8'sb00010000, 8'sb00010011, 8'sb00001011, 8'sb00001010, 8'sb00001001, 8'sb00001011, 8'sb00000011, 8'sb11110101, 8'sb00000011, 8'sb00001011, 8'sb00001001, 8'sb00000111, 8'sb11110111, 8'sb11111111, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00011110, 8'sb00100011, 8'sb00011010, 8'sb00010101, 8'sb00110000, 8'sb00101101, 8'sb00010001, 8'sb00100001, 8'sb00100101, 8'sb00010000, 8'sb00001100, 8'sb00010000, 8'sb00010001, 8'sb00010010, 8'sb00100010, 8'sb00100111, 8'sb00100000, 8'sb00011011, 8'sb00100100, 8'sb00011110, 8'sb00011001, 8'sb00010011, 8'sb00010101, 8'sb00001001, 8'sb00010010, 8'sb00010011, 8'sb00010011, 8'sb00010010, 8'sb00011010, 8'sb00011100, 8'sb00001001, 8'sb00010100, 8'sb00011011, 8'sb00100010, 8'sb00010111, 8'sb00001110, 8'sb00001101, 8'sb00001001, 8'sb00001110, 8'sb00010010, 8'sb00010011, 8'sb00001111, 8'sb00000101, 8'sb00001000, 8'sb00011100, 8'sb00011110, 8'sb00100100, 8'sb00101011, 8'sb00011011, 8'sb00010010, 8'sb00001011, 8'sb00000111, 8'sb00010101, 8'sb00010100, 8'sb00010000, 8'sb00010001, 8'sb00000010, 8'sb11101010, 8'sb11101111, 8'sb00000001, 8'sb00001000, 8'sb00000111, 8'sb00000110, 8'sb00001100, 8'sb00000000, 8'sb00001000, 8'sb00010010, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00001100, 8'sb00000000, 8'sb11110111, 8'sb11100101, 8'sb11100100, 8'sb11101101, 8'sb11101111, 8'sb11111100, 8'sb00000110, 8'sb00001111, 8'sb00010011, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00001111, 8'sb00001001, 8'sb11111111, 8'sb11111100, 8'sb00010000, 8'sb00010000, 8'sb00011110, 8'sb00010100, 8'sb00010011, 8'sb00010011, 8'sb00010010, 8'sb00010100, 8'sb00010001, 8'sb00010010, 8'sb00001101, 8'sb00001110, 8'sb00010100, 8'sb00010101, 8'sb00010000, 8'sb00001110, 8'sb00010011, 8'sb00010010, 8'sb00010001, 8'sb00010000,
    8'sb00001100, 8'sb00001101, 8'sb00001101, 8'sb00001101, 8'sb00001011, 8'sb00001011, 8'sb00001110, 8'sb00001100, 8'sb00001010, 8'sb00001011, 8'sb00001100, 8'sb00001011, 8'sb00001111, 8'sb00001111, 8'sb00001101, 8'sb00001111, 8'sb00001110, 8'sb00001101, 8'sb00001111, 8'sb00010110, 8'sb00011010, 8'sb00010011, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00001110, 8'sb00001101, 8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00001111, 8'sb00010100, 8'sb00011000, 8'sb00011110, 8'sb00011000, 8'sb00000010, 8'sb00001111, 8'sb00010111, 8'sb00010101, 8'sb00001111, 8'sb00010011, 8'sb00001101, 8'sb00001110, 8'sb00001011, 8'sb00010000, 8'sb00010010, 8'sb00011111, 8'sb00001100, 8'sb00001100, 8'sb00010111, 8'sb00010010, 8'sb00000100, 8'sb00000111, 8'sb00001101, 8'sb00010011, 8'sb00001011, 8'sb00001100, 8'sb00001010, 8'sb00000101, 8'sb00001010, 8'sb00001111, 8'sb00010000, 8'sb00000111, 8'sb00000000, 8'sb11111111, 8'sb00000001, 8'sb00000100, 8'sb00000111, 8'sb00000110, 8'sb00001111, 8'sb00001011, 8'sb00000111, 8'sb00001000, 8'sb00010100, 8'sb00100010, 8'sb00010100, 8'sb11110000, 8'sb11101110, 8'sb00000001, 8'sb00000100, 8'sb00000010, 8'sb11111101, 8'sb00000010, 8'sb00001110, 8'sb00001011, 8'sb00001010, 8'sb00000110, 8'sb00000100, 8'sb00010100, 8'sb00101011, 8'sb00011010, 8'sb00001100, 8'sb00010010, 8'sb00010100, 8'sb00010000, 8'sb00001000, 8'sb00001111, 8'sb00001111, 8'sb00001111, 8'sb00001111, 8'sb00000110, 8'sb00001111, 8'sb00010000, 8'sb00011110, 8'sb00100010, 8'sb00010011, 8'sb00011001, 8'sb00001011, 8'sb00001001, 8'sb00001100, 8'sb00001110, 8'sb00001110, 8'sb00001100, 8'sb00001110, 8'sb00001100, 8'sb00000110, 8'sb00010011, 8'sb00011010, 8'sb00101011, 8'sb00010110, 8'sb00011011, 8'sb00011101, 8'sb00011000, 8'sb00011000, 8'sb00010110, 8'sb00010000, 8'sb00001111, 8'sb00010011, 8'sb00011011, 8'sb00010011, 8'sb11111111, 8'sb00001100, 8'sb00001111, 8'sb00001011, 8'sb00010001, 8'sb00010000, 8'sb00011000, 8'sb00010111, 8'sb00011000, 8'sb00001110, 8'sb00001011, 8'sb00010011, 8'sb00011000, 8'sb00001101, 8'sb00001010, 8'sb11111101, 8'sb00010100, 8'sb00011100, 8'sb00010001, 8'sb00011001, 8'sb00011000, 8'sb00011111, 8'sb00001111, 8'sb00001111, 8'sb00001101, 8'sb00010001, 8'sb00010110, 8'sb00001100, 8'sb00010110, 8'sb00010010, 8'sb00001000, 8'sb00001101, 8'sb00010101, 8'sb00101001, 8'sb00100011, 8'sb00010111, 8'sb00010000, 8'sb00001101, 8'sb00001100, 8'sb00001111, 8'sb00001101, 8'sb00001001, 8'sb00001100, 8'sb00010011, 8'sb00010010, 8'sb00010100, 8'sb00001110, 8'sb00010100, 8'sb00010101, 8'sb00010011, 8'sb00001111, 8'sb00001110, 8'sb00001100, 8'sb00001011, 8'sb00001110, 8'sb00001101, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00001101, 8'sb00000110, 8'sb00000101, 8'sb00001101, 8'sb00001110, 8'sb00001111, 8'sb00001100,
    8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00001101, 8'sb00001101, 8'sb00010001, 8'sb00001101, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00001101, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00010000, 8'sb00001110, 8'sb00001100, 8'sb00010001, 8'sb00001110, 8'sb00000111, 8'sb00001010, 8'sb00001001, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00001111, 8'sb00001101, 8'sb00001101, 8'sb00001101, 8'sb00001100, 8'sb11111111, 8'sb11111100, 8'sb00000001, 8'sb00000011, 8'sb00010100, 8'sb00011110, 8'sb00010100, 8'sb00010001, 8'sb00001111, 8'sb00001101, 8'sb00001011, 8'sb00010011, 8'sb00011010, 8'sb00100000, 8'sb00010100, 8'sb11111111, 8'sb11110011, 8'sb00000101, 8'sb00001001, 8'sb00011101, 8'sb00100011, 8'sb00010000, 8'sb00001111, 8'sb00001101, 8'sb00001111, 8'sb00001101, 8'sb00010001, 8'sb00010110, 8'sb00101110, 8'sb00000000, 8'sb11100100, 8'sb11110100, 8'sb00000110, 8'sb00001010, 8'sb00100110, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00010100, 8'sb00010101, 8'sb00010010, 8'sb00100010, 8'sb00101010, 8'sb00000001, 8'sb11101110, 8'sb11111000, 8'sb00000011, 8'sb00010110, 8'sb00010010, 8'sb00001100, 8'sb00001100, 8'sb00001111, 8'sb00011000, 8'sb00010001, 8'sb00001110, 8'sb00100011, 8'sb00100001, 8'sb00010010, 8'sb00001010, 8'sb00001101, 8'sb00000110, 8'sb00001100, 8'sb00001101, 8'sb00001110, 8'sb00001110, 8'sb00001000, 8'sb00000111, 8'sb00001110, 8'sb00011100, 8'sb00011100, 8'sb00100101, 8'sb00000100, 8'sb00001100, 8'sb00001001, 8'sb00001000, 8'sb00010000, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00000010, 8'sb00001010, 8'sb00010011, 8'sb00010101, 8'sb00100101, 8'sb00011011, 8'sb00001101, 8'sb00001001, 8'sb00010000, 8'sb00010001, 8'sb00010011, 8'sb00001101, 8'sb00010000, 8'sb00001101, 8'sb00001111, 8'sb00010001, 8'sb00011000, 8'sb00010100, 8'sb00001110, 8'sb00010010, 8'sb00001110, 8'sb00001110, 8'sb00010100, 8'sb00011000, 8'sb00001101, 8'sb00010000, 8'sb00010001, 8'sb00001001, 8'sb00001000, 8'sb00010011, 8'sb00010100, 8'sb00001011, 8'sb00000100, 8'sb00010101, 8'sb00010100, 8'sb00010100, 8'sb00010010, 8'sb00010001, 8'sb00001011, 8'sb00001100, 8'sb00010001, 8'sb00001011, 8'sb00001100, 8'sb00010100, 8'sb00010001, 8'sb00001010, 8'sb00001110, 8'sb00001001, 8'sb00010111, 8'sb00010000, 8'sb00001111, 8'sb00001101, 8'sb00001100, 8'sb00010000, 8'sb00010000, 8'sb00001110, 8'sb00000101, 8'sb11111111, 8'sb00000101, 8'sb00001000, 8'sb00001001, 8'sb00001110, 8'sb00010011, 8'sb00011010, 8'sb00001100, 8'sb00010000, 8'sb00010000, 8'sb00001110, 8'sb00001111, 8'sb00001110, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00000111, 8'sb00000001, 8'sb00000011, 8'sb00001001, 8'sb00001010, 8'sb00001111, 8'sb00001110, 8'sb00001101, 8'sb00001101,
    8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00010000, 8'sb00001101, 8'sb00010000, 8'sb00010001, 8'sb00001110, 8'sb00001101, 8'sb00001111, 8'sb00001110, 8'sb00010000, 8'sb00010001, 8'sb00010001, 8'sb00001110, 8'sb00001100, 8'sb00001101, 8'sb00001011, 8'sb00001111, 8'sb00001100, 8'sb00001101, 8'sb00010000, 8'sb00001111, 8'sb00010001, 8'sb00010000, 8'sb00001100, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00001001, 8'sb00000010, 8'sb00000001, 8'sb00010010, 8'sb00000111, 8'sb00001001, 8'sb00000100, 8'sb00001011, 8'sb00001101, 8'sb00001101, 8'sb00010001, 8'sb00010011, 8'sb00011101, 8'sb00011011, 8'sb00011000, 8'sb00011001, 8'sb00001101, 8'sb00011011, 8'sb00010011, 8'sb00010011, 8'sb00010101, 8'sb00000111, 8'sb00000111, 8'sb00001110, 8'sb00001110, 8'sb00010100, 8'sb00011101, 8'sb00011001, 8'sb00010111, 8'sb00011000, 8'sb00000110, 8'sb00101011, 8'sb00010001, 8'sb00011100, 8'sb00010101, 8'sb00001101, 8'sb00000111, 8'sb00001100, 8'sb00010010, 8'sb00011101, 8'sb00010011, 8'sb00000001, 8'sb00000011, 8'sb00001011, 8'sb00000110, 8'sb00111111, 8'sb00110111, 8'sb00100110, 8'sb00011101, 8'sb00001100, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00010101, 8'sb00000100, 8'sb00000011, 8'sb11111110, 8'sb11110110, 8'sb11101110, 8'sb00000101, 8'sb00001011, 8'sb00001001, 8'sb00001100, 8'sb00010011, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00001001, 8'sb00000000, 8'sb00000100, 8'sb11111110, 8'sb11111100, 8'sb11111101, 8'sb00000000, 8'sb00010011, 8'sb00100001, 8'sb00100001, 8'sb00001111, 8'sb00001111, 8'sb00001100, 8'sb00010001, 8'sb00001101, 8'sb00000011, 8'sb00001011, 8'sb00000000, 8'sb11111010, 8'sb00000110, 8'sb00001010, 8'sb00010001, 8'sb00011001, 8'sb00010111, 8'sb00001110, 8'sb00001110, 8'sb00010001, 8'sb00010110, 8'sb00001111, 8'sb00000001, 8'sb00001100, 8'sb00000111, 8'sb00000011, 8'sb00001100, 8'sb00001010, 8'sb00001100, 8'sb00001001, 8'sb00001011, 8'sb00001100, 8'sb00001101, 8'sb00001100, 8'sb00010100, 8'sb00010111, 8'sb00011001, 8'sb00011110, 8'sb00011000, 8'sb00100011, 8'sb00011000, 8'sb00001100, 8'sb00000000, 8'sb00000001, 8'sb11111111, 8'sb00001101, 8'sb00010001, 8'sb00001101, 8'sb00010000, 8'sb00011010, 8'sb00100101, 8'sb00010100, 8'sb00001110, 8'sb00001110, 8'sb00011000, 8'sb00010100, 8'sb00010000, 8'sb11111110, 8'sb00000011, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00001110, 8'sb00010010, 8'sb00011000, 8'sb00010100, 8'sb00010010, 8'sb00010000, 8'sb00000110, 8'sb00001011, 8'sb00000111, 8'sb00000001, 8'sb00001000, 8'sb00010000, 8'sb00001110, 8'sb00001110, 8'sb00010001, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00001100, 8'sb00001101, 8'sb00010110, 8'sb00010100, 8'sb00010110, 8'sb00001110, 8'sb00010000, 8'sb00010000, 8'sb00001110,
    8'sb00010011, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00010011, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010100, 8'sb00010100, 8'sb00010001, 8'sb00001001, 8'sb00001010, 8'sb00001000, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00010011, 8'sb00010001, 8'sb00001111, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00001110, 8'sb00001101, 8'sb00000100, 8'sb00000111, 8'sb00001110, 8'sb00001100, 8'sb00010011, 8'sb00010010, 8'sb00010010, 8'sb00001110, 8'sb00010010, 8'sb00010010, 8'sb00010101, 8'sb00011011, 8'sb00010011, 8'sb00001100, 8'sb00000110, 8'sb00010011, 8'sb00010000, 8'sb00001110, 8'sb00010101, 8'sb00010011, 8'sb00010001, 8'sb00010010, 8'sb00010001, 8'sb00010000, 8'sb00010111, 8'sb00100000, 8'sb00011111, 8'sb00100000, 8'sb00010101, 8'sb00010101, 8'sb00010010, 8'sb00010010, 8'sb00010101, 8'sb00010010, 8'sb00010000, 8'sb00010001, 8'sb00001010, 8'sb00001111, 8'sb00010010, 8'sb00001100, 8'sb00010011, 8'sb00001111, 8'sb00001000, 8'sb00000101, 8'sb11111100, 8'sb11111110, 8'sb00010011, 8'sb00010100, 8'sb00010011, 8'sb00001111, 8'sb11111101, 8'sb11110001, 8'sb11101110, 8'sb11100100, 8'sb11100010, 8'sb11110101, 8'sb11111010, 8'sb11110111, 8'sb11111100, 8'sb00000000, 8'sb00001110, 8'sb00010010, 8'sb00001111, 8'sb00010000, 8'sb11110111, 8'sb11100001, 8'sb11110110, 8'sb00000011, 8'sb00010001, 8'sb00001010, 8'sb00000101, 8'sb00000111, 8'sb00010000, 8'sb00000111, 8'sb00010011, 8'sb00011001, 8'sb00010011, 8'sb00001011, 8'sb00000010, 8'sb00010000, 8'sb00011010, 8'sb00010011, 8'sb00011001, 8'sb00010101, 8'sb00001011, 8'sb00000011, 8'sb00010100, 8'sb00001110, 8'sb00011010, 8'sb00011000, 8'sb00010011, 8'sb00001101, 8'sb00010000, 8'sb00010100, 8'sb00011011, 8'sb00010101, 8'sb00011000, 8'sb00011011, 8'sb00001111, 8'sb00000111, 8'sb00000010, 8'sb00001000, 8'sb00011100, 8'sb00010101, 8'sb00001111, 8'sb00010001, 8'sb00010000, 8'sb00001100, 8'sb00010010, 8'sb00010100, 8'sb00010101, 8'sb00010110, 8'sb00001110, 8'sb00001111, 8'sb00000100, 8'sb00010100, 8'sb00011010, 8'sb00010011, 8'sb00010010, 8'sb00001111, 8'sb00001100, 8'sb00010010, 8'sb00010010, 8'sb00010010, 8'sb00010010, 8'sb00010100, 8'sb00001010, 8'sb00010001, 8'sb00010111, 8'sb00011011, 8'sb00010011, 8'sb00010000, 8'sb00010011, 8'sb00001111, 8'sb00001100, 8'sb00001000, 8'sb00001001, 8'sb00001100, 8'sb00001000, 8'sb00001100, 8'sb00010001, 8'sb00010100, 8'sb00010001, 8'sb00010001, 8'sb00010001, 8'sb00010001, 8'sb00001111, 8'sb00010010, 8'sb00010011, 8'sb00010001, 8'sb00010001, 8'sb00010110, 8'sb00010000, 8'sb00010110, 8'sb00010011, 8'sb00010000, 8'sb00010000, 8'sb00010000, 8'sb00010011, 8'sb00001111,
    8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00010010, 8'sb00001111, 8'sb00010001, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00010001, 8'sb00010001, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00001101, 8'sb00001110, 8'sb00001111, 8'sb00010001, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00010100, 8'sb00010011, 8'sb00000110, 8'sb11111100, 8'sb11110100, 8'sb11110001, 8'sb11111001, 8'sb00000011, 8'sb00001011, 8'sb00010001, 8'sb00010000, 8'sb00001110, 8'sb00010100, 8'sb00011000, 8'sb00010101, 8'sb00011011, 8'sb00010001, 8'sb00011111, 8'sb00010001, 8'sb00010100, 8'sb00001100, 8'sb00001101, 8'sb00000101, 8'sb00001100, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00010100, 8'sb00010010, 8'sb00010100, 8'sb00011001, 8'sb00011011, 8'sb00010101, 8'sb00010010, 8'sb00011000, 8'sb00010001, 8'sb00011000, 8'sb00001010, 8'sb00010001, 8'sb00001111, 8'sb00011001, 8'sb00010001, 8'sb00001111, 8'sb00010010, 8'sb00010100, 8'sb00001111, 8'sb00010100, 8'sb00010101, 8'sb00011101, 8'sb00100011, 8'sb00010001, 8'sb00001001, 8'sb00010001, 8'sb00010011, 8'sb00010100, 8'sb00010000, 8'sb00010001, 8'sb00000101, 8'sb00001011, 8'sb00001101, 8'sb00100110, 8'sb00100000, 8'sb00010011, 8'sb00001101, 8'sb00001010, 8'sb00001010, 8'sb00010010, 8'sb00001111, 8'sb00010011, 8'sb00001001, 8'sb00000111, 8'sb00001010, 8'sb00001010, 8'sb00001110, 8'sb00010111, 8'sb00010110, 8'sb00011011, 8'sb00010101, 8'sb00001011, 8'sb00010000, 8'sb00010001, 8'sb00010000, 8'sb00010100, 8'sb00010001, 8'sb00001100, 8'sb00010000, 8'sb00001001, 8'sb00001000, 8'sb00001010, 8'sb00010100, 8'sb00010001, 8'sb00011000, 8'sb00010011, 8'sb00001110, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00001101, 8'sb11110011, 8'sb11110110, 8'sb11111010, 8'sb11111000, 8'sb00000010, 8'sb00000100, 8'sb00000110, 8'sb00010000, 8'sb00001000, 8'sb00001011, 8'sb00001110, 8'sb00010001, 8'sb00010011, 8'sb00000101, 8'sb11110011, 8'sb11111001, 8'sb11111010, 8'sb11111011, 8'sb11111101, 8'sb11111111, 8'sb00000100, 8'sb00001000, 8'sb11111110, 8'sb00001100, 8'sb00010010, 8'sb00010010, 8'sb00010011, 8'sb00010100, 8'sb00010010, 8'sb00001000, 8'sb00000111, 8'sb11111101, 8'sb00000010, 8'sb11111100, 8'sb11110110, 8'sb11111010, 8'sb00000010, 8'sb00001101, 8'sb00001110, 8'sb00010000, 8'sb00010001, 8'sb00011111, 8'sb00100101, 8'sb00010111, 8'sb00011010, 8'sb00011000, 8'sb00010000, 8'sb00010000, 8'sb00000100, 8'sb00001101, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00010001, 8'sb00010010, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00010100, 8'sb00011000, 8'sb00011000, 8'sb00010110, 8'sb00010010, 8'sb00010010, 8'sb00001110, 8'sb00010001,
    8'sb00001010, 8'sb00001100, 8'sb00001101, 8'sb00001000, 8'sb00001010, 8'sb00001001, 8'sb00001011, 8'sb00001011, 8'sb00001010, 8'sb00001101, 8'sb00001100, 8'sb00001010, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00001000, 8'sb00001011, 8'sb00001000, 8'sb00001111, 8'sb00010101, 8'sb00011010, 8'sb00010011, 8'sb00010111, 8'sb00010001, 8'sb00001010, 8'sb00001110, 8'sb00001011, 8'sb00001100, 8'sb00001001, 8'sb00001010, 8'sb00000111, 8'sb00000111, 8'sb00010011, 8'sb00010001, 8'sb00000111, 8'sb00000100, 8'sb00001001, 8'sb00000011, 8'sb00001001, 8'sb00001111, 8'sb00001100, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00000101, 8'sb00010000, 8'sb00001110, 8'sb00001000, 8'sb00001111, 8'sb00001001, 8'sb00001001, 8'sb00001101, 8'sb00000100, 8'sb00001001, 8'sb00000111, 8'sb00001001, 8'sb00001010, 8'sb00001101, 8'sb00001101, 8'sb00010001, 8'sb00001001, 8'sb00010001, 8'sb00011001, 8'sb00011010, 8'sb00011010, 8'sb00001101, 8'sb00001100, 8'sb00001001, 8'sb11111101, 8'sb00001001, 8'sb00001100, 8'sb00010001, 8'sb00011111, 8'sb00011001, 8'sb00001001, 8'sb00001011, 8'sb11111111, 8'sb11111010, 8'sb00001011, 8'sb00001100, 8'sb00010011, 8'sb00011001, 8'sb00001101, 8'sb00001100, 8'sb00001001, 8'sb00010100, 8'sb00100100, 8'sb00100000, 8'sb00001000, 8'sb00001000, 8'sb11111010, 8'sb11101100, 8'sb11111110, 8'sb00000101, 8'sb00011111, 8'sb00101110, 8'sb00011100, 8'sb00001001, 8'sb00001101, 8'sb00001101, 8'sb00011111, 8'sb00110111, 8'sb00101100, 8'sb00010010, 8'sb11101111, 8'sb00000001, 8'sb00011101, 8'sb00100010, 8'sb00011011, 8'sb00010111, 8'sb00010011, 8'sb00001010, 8'sb00001010, 8'sb00001010, 8'sb00010011, 8'sb00100010, 8'sb00111111, 8'sb00111010, 8'sb00001111, 8'sb00011100, 8'sb00011101, 8'sb00010010, 8'sb00001110, 8'sb00000101, 8'sb00010010, 8'sb00001101, 8'sb00001100, 8'sb00000011, 8'sb00000101, 8'sb11111111, 8'sb00000111, 8'sb00101001, 8'sb00110010, 8'sb00010111, 8'sb00001000, 8'sb00010010, 8'sb00000110, 8'sb00001101, 8'sb00010110, 8'sb00001011, 8'sb00001010, 8'sb00001001, 8'sb00000111, 8'sb00000110, 8'sb00000010, 8'sb00001010, 8'sb00010100, 8'sb00011001, 8'sb00010010, 8'sb00001010, 8'sb00001101, 8'sb00011101, 8'sb00010100, 8'sb00001010, 8'sb00001010, 8'sb00001011, 8'sb00000111, 8'sb00001111, 8'sb00010010, 8'sb00001101, 8'sb00001011, 8'sb00000110, 8'sb00000101, 8'sb00010101, 8'sb00011010, 8'sb00011011, 8'sb00010000, 8'sb00001100, 8'sb00001001, 8'sb00001011, 8'sb00001011, 8'sb00000110, 8'sb00000011, 8'sb00000111, 8'sb00001011, 8'sb00010010, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00001100, 8'sb00001001, 8'sb00001100, 8'sb00001010, 8'sb00001010, 8'sb00001001, 8'sb00001011, 8'sb00001010, 8'sb00001101, 8'sb00010011, 8'sb00010010, 8'sb00001101, 8'sb00001111, 8'sb00001101, 8'sb00001100, 8'sb00001000, 8'sb00001100,
    8'sb00001101, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00001111, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00000100, 8'sb11111111, 8'sb00000001, 8'sb00000100, 8'sb00000011, 8'sb00000111, 8'sb00000111, 8'sb00001010, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00010010, 8'sb00010011, 8'sb00010100, 8'sb00001101, 8'sb00001110, 8'sb00010111, 8'sb00010110, 8'sb00001100, 8'sb00001010, 8'sb00001001, 8'sb00001100, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00010110, 8'sb00010000, 8'sb00010101, 8'sb00010100, 8'sb00001110, 8'sb00001000, 8'sb00000100, 8'sb11111110, 8'sb00001001, 8'sb00010101, 8'sb00010001, 8'sb00001110, 8'sb00010001, 8'sb00001110, 8'sb00011000, 8'sb00010111, 8'sb00001111, 8'sb00001100, 8'sb00001110, 8'sb00001100, 8'sb00010000, 8'sb00100000, 8'sb00011001, 8'sb00100100, 8'sb00011011, 8'sb00010001, 8'sb00001110, 8'sb00010001, 8'sb00010001, 8'sb00010001, 8'sb00010000, 8'sb00011100, 8'sb00011100, 8'sb00110000, 8'sb00100101, 8'sb00011010, 8'sb00011011, 8'sb00010100, 8'sb00011000, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00001100, 8'sb00010111, 8'sb00010101, 8'sb00011100, 8'sb00011110, 8'sb00011010, 8'sb00010011, 8'sb00010011, 8'sb00000000, 8'sb00010000, 8'sb00010100, 8'sb00010001, 8'sb00010001, 8'sb00001100, 8'sb11111000, 8'sb00001011, 8'sb00010001, 8'sb00010101, 8'sb00011111, 8'sb00101000, 8'sb00010011, 8'sb00000011, 8'sb00000110, 8'sb00001001, 8'sb00010000, 8'sb00001111, 8'sb00011000, 8'sb00010100, 8'sb00000100, 8'sb00000010, 8'sb11111100, 8'sb00100001, 8'sb00101101, 8'sb00010000, 8'sb11111010, 8'sb00000101, 8'sb00010101, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00011000, 8'sb00011000, 8'sb00010001, 8'sb00000110, 8'sb00000010, 8'sb00000110, 8'sb11111001, 8'sb11101110, 8'sb11111110, 8'sb00000001, 8'sb00001000, 8'sb00001000, 8'sb00001101, 8'sb00001101, 8'sb00010010, 8'sb00001101, 8'sb00010000, 8'sb00000111, 8'sb00000110, 8'sb00000000, 8'sb00000011, 8'sb00001001, 8'sb00000110, 8'sb00000010, 8'sb00000010, 8'sb00001000, 8'sb00001110, 8'sb00010010, 8'sb00010010, 8'sb00001100, 8'sb00010000, 8'sb00001010, 8'sb00000110, 8'sb00001111, 8'sb00010011, 8'sb00010100, 8'sb00011100, 8'sb00010101, 8'sb00010010, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00010001, 8'sb00010101, 8'sb00010110, 8'sb00000110, 8'sb00001111, 8'sb00001110, 8'sb00010001, 8'sb00010001, 8'sb00010001, 8'sb00001111, 8'sb00001101, 8'sb00001101, 8'sb00010001, 8'sb00001101, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00001100, 8'sb00001111, 8'sb00001100, 8'sb00001111, 8'sb00010001, 8'sb00010001, 8'sb00001101,
    8'sb00010011, 8'sb00010110, 8'sb00010101, 8'sb00010010, 8'sb00010101, 8'sb00010101, 8'sb00010011, 8'sb00010100, 8'sb00010010, 8'sb00010010, 8'sb00010011, 8'sb00010011, 8'sb00010100, 8'sb00010101, 8'sb00010110, 8'sb00010100, 8'sb00010101, 8'sb00010101, 8'sb00010001, 8'sb00001000, 8'sb00000101, 8'sb00001001, 8'sb00001010, 8'sb00001111, 8'sb00010011, 8'sb00010101, 8'sb00010010, 8'sb00010101, 8'sb00010100, 8'sb00010011, 8'sb00010011, 8'sb00010000, 8'sb00000001, 8'sb11111010, 8'sb11111101, 8'sb00000110, 8'sb00000011, 8'sb00001001, 8'sb00010010, 8'sb00011010, 8'sb00001111, 8'sb00010100, 8'sb00010011, 8'sb00010100, 8'sb00010010, 8'sb00000011, 8'sb11110111, 8'sb00000001, 8'sb00001110, 8'sb00000110, 8'sb00001000, 8'sb00010000, 8'sb00001011, 8'sb00010011, 8'sb00010101, 8'sb00010100, 8'sb00010101, 8'sb00010001, 8'sb00001110, 8'sb00000011, 8'sb11111110, 8'sb11111111, 8'sb00010110, 8'sb00011011, 8'sb00010111, 8'sb00010001, 8'sb00010000, 8'sb00001111, 8'sb00100101, 8'sb00010101, 8'sb00010010, 8'sb00010011, 8'sb00001110, 8'sb00000111, 8'sb00000111, 8'sb00001010, 8'sb00011000, 8'sb00100001, 8'sb00001011, 8'sb00000000, 8'sb00001100, 8'sb00011110, 8'sb00101101, 8'sb00010111, 8'sb00010011, 8'sb00010011, 8'sb00010110, 8'sb00010011, 8'sb00001100, 8'sb00001011, 8'sb00011000, 8'sb00010100, 8'sb00000110, 8'sb11100000, 8'sb11011101, 8'sb11101100, 8'sb00001000, 8'sb00010110, 8'sb00010101, 8'sb00010110, 8'sb00010011, 8'sb00001101, 8'sb00010010, 8'sb00001110, 8'sb00001100, 8'sb00001101, 8'sb00010000, 8'sb00001101, 8'sb11110100, 8'sb11111000, 8'sb00001101, 8'sb00010001, 8'sb00010101, 8'sb00010001, 8'sb00010010, 8'sb00001011, 8'sb00000100, 8'sb00001001, 8'sb00001101, 8'sb00010111, 8'sb00001101, 8'sb00001111, 8'sb11111001, 8'sb00000000, 8'sb00001001, 8'sb00010011, 8'sb00010110, 8'sb00010001, 8'sb00010011, 8'sb00010101, 8'sb00000111, 8'sb00001000, 8'sb00010111, 8'sb00001111, 8'sb00001100, 8'sb00010000, 8'sb11111111, 8'sb00000011, 8'sb00001101, 8'sb00010100, 8'sb00010101, 8'sb00001110, 8'sb00000100, 8'sb00001000, 8'sb00010010, 8'sb00001111, 8'sb00001001, 8'sb00001111, 8'sb00010001, 8'sb00010001, 8'sb00000100, 8'sb00001010, 8'sb00010011, 8'sb00010110, 8'sb00010101, 8'sb00010011, 8'sb00010011, 8'sb00001001, 8'sb00010011, 8'sb00001111, 8'sb00001001, 8'sb00000111, 8'sb00010101, 8'sb00011000, 8'sb00001100, 8'sb00010001, 8'sb00010010, 8'sb00010101, 8'sb00010100, 8'sb00010011, 8'sb00001110, 8'sb00001011, 8'sb00001000, 8'sb00001100, 8'sb00001010, 8'sb00000101, 8'sb00001000, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00010011, 8'sb00010010, 8'sb00010100, 8'sb00010010, 8'sb00010101, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00001100, 8'sb00010001, 8'sb00010001, 8'sb00010110, 8'sb00010110, 8'sb00010100,
    8'sb00001101, 8'sb00001011, 8'sb00001101, 8'sb00001111, 8'sb00001011, 8'sb00001111, 8'sb00001100, 8'sb00001101, 8'sb00001111, 8'sb00001101, 8'sb00001011, 8'sb00001011, 8'sb00001100, 8'sb00001011, 8'sb00001010, 8'sb00001010, 8'sb00001111, 8'sb00001110, 8'sb00010011, 8'sb00011011, 8'sb00011111, 8'sb00011111, 8'sb00011010, 8'sb00010011, 8'sb00001101, 8'sb00001101, 8'sb00001101, 8'sb00001010, 8'sb00001110, 8'sb00001101, 8'sb00001101, 8'sb00010100, 8'sb00011100, 8'sb00011011, 8'sb00011000, 8'sb00010111, 8'sb00010110, 8'sb00001101, 8'sb00000110, 8'sb00000111, 8'sb00001110, 8'sb00001111, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00010000, 8'sb00010111, 8'sb00001011, 8'sb00001110, 8'sb00001001, 8'sb00000101, 8'sb00001000, 8'sb00000101, 8'sb00001000, 8'sb00010001, 8'sb00001110, 8'sb00001110, 8'sb00001001, 8'sb00000011, 8'sb00010001, 8'sb00010100, 8'sb00001011, 8'sb00000011, 8'sb00010001, 8'sb00001001, 8'sb00000111, 8'sb00010010, 8'sb00010000, 8'sb00011000, 8'sb00001101, 8'sb00001011, 8'sb00001000, 8'sb00001011, 8'sb00010001, 8'sb00000100, 8'sb00001100, 8'sb00010111, 8'sb00001100, 8'sb00000111, 8'sb00000000, 8'sb00001001, 8'sb00001010, 8'sb00010110, 8'sb00001100, 8'sb00001110, 8'sb00001011, 8'sb00000010, 8'sb11110111, 8'sb11111111, 8'sb00011000, 8'sb00010010, 8'sb11111111, 8'sb00000010, 8'sb00000111, 8'sb00000111, 8'sb00010000, 8'sb00010110, 8'sb00001011, 8'sb00001100, 8'sb00001100, 8'sb00001001, 8'sb00001000, 8'sb00001110, 8'sb00010010, 8'sb00001011, 8'sb00001110, 8'sb00000011, 8'sb00001110, 8'sb00010010, 8'sb00011010, 8'sb00100001, 8'sb00001110, 8'sb00001110, 8'sb00010001, 8'sb00011010, 8'sb00010111, 8'sb00000011, 8'sb00001001, 8'sb11111101, 8'sb00000110, 8'sb00001010, 8'sb00010011, 8'sb00001110, 8'sb00101010, 8'sb00100110, 8'sb00001110, 8'sb00001100, 8'sb00001110, 8'sb00011010, 8'sb00101001, 8'sb00101000, 8'sb00101010, 8'sb00010011, 8'sb00001100, 8'sb00010100, 8'sb00010110, 8'sb00010001, 8'sb00101100, 8'sb00011101, 8'sb00001110, 8'sb00001011, 8'sb00010000, 8'sb00011010, 8'sb00011010, 8'sb00101000, 8'sb00101111, 8'sb00100010, 8'sb00010110, 8'sb00010010, 8'sb00011000, 8'sb00010100, 8'sb00011100, 8'sb00010010, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00001010, 8'sb00000001, 8'sb00001001, 8'sb00010000, 8'sb00011010, 8'sb00010110, 8'sb00010011, 8'sb00010011, 8'sb00011001, 8'sb00010000, 8'sb00001111, 8'sb00001100, 8'sb00001110, 8'sb00001101, 8'sb00000111, 8'sb00000011, 8'sb00000000, 8'sb00000010, 8'sb00000010, 8'sb00001010, 8'sb00001011, 8'sb00001011, 8'sb00000101, 8'sb00001100, 8'sb00001100, 8'sb00001011, 8'sb00001010, 8'sb00001010, 8'sb00001011, 8'sb00001101, 8'sb00001010, 8'sb00001001, 8'sb00001010, 8'sb00001000, 8'sb00001001, 8'sb00001100, 8'sb00001001, 8'sb00001100, 8'sb00001010, 8'sb00001100
    };

    localparam signed [8*30-1:0] biases_HL_param = {
    8'sb00010100, 8'sb00010011, 8'sb00010000, 8'sb00001010, 8'sb00010010, 8'sb00000011, 8'sb00000010, 8'sb00001000, 8'sb00010001, 8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00010010, 8'sb00000100, 8'sb00011000, 8'sb00010100, 8'sb00001010, 8'sb00001111, 8'sb00010100, 8'sb00000101, 8'sb00000111, 8'sb00010010, 8'sb00001110, 8'sb00001111, 8'sb00001001, 8'sb00001001, 8'sb00010111, 8'sb00001011, 8'sb00000000, 8'sb00010010
    };

    integer i, j;

    // Assign values to weights and biases
    always @(*) begin
        // Assign weights from the flattened localparam to the output
        for (i = 0; i < 30; i = i + 1) begin
            for (j = 0; j < 196; j = j + 1) begin
                weights_HL[(i * 196 + j) * 8] = weights_HL_param[(i * 196 + j)*8];
                weights_HL[(i * 196 + j) * 8 + 1] = weights_HL_param[(i * 196 + j)*8 + 1];
                weights_HL[(i * 196 + j) * 8 + 2] = weights_HL_param[(i * 196 + j)*8 + 2];
                weights_HL[(i * 196 + j) * 8 + 3] = weights_HL_param[(i * 196 + j)*8 + 3];
                weights_HL[(i * 196 + j) * 8 + 4] = weights_HL_param[(i * 196 + j)*8 + 4];
                weights_HL[(i * 196 + j) * 8 + 5] = weights_HL_param[(i * 196 + j)*8 + 5];
                weights_HL[(i * 196 + j) * 8 + 6] = weights_HL_param[(i * 196 + j)*8 + 6];
                weights_HL[(i * 196 + j) * 8 + 7] = weights_HL_param[(i * 196 + j)*8 + 7];
            end
            biases_HL[i * 8] = biases_HL_param[i * 8];
            biases_HL[i * 8 + 1] = biases_HL_param[i * 8 + 1];
            biases_HL[i * 8 + 2] = biases_HL_param[i * 8 + 2];
            biases_HL[i * 8 + 3] = biases_HL_param[i * 8 + 3];
            biases_HL[i * 8 + 4] = biases_HL_param[i * 8 + 4];
            biases_HL[i * 8 + 5] = biases_HL_param[i * 8 + 5];
            biases_HL[i * 8 + 6] = biases_HL_param[i * 8 + 6];
            biases_HL[i * 8 + 7] = biases_HL_param[i * 8 + 7];
        end
    end

endmodule
