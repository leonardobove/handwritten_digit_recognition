//////////////////////////////////////////////////////////////////////////////////

/**********
* 1st dense layer implementation (hidden layer)
*
* Inputs: clk => clock signal, enable => enable signal, 
*         reset => active high sync reset, pooled_img => in vector, 
*
* Outputs: hidden_out => dense layer output
*          layer_done => done signal
* 
***********/


module hidden_layer #(
    parameter averaged_pixels_nr = 196,
    parameter WIDTH = 8,
    parameter HL_neurons = 32
	)(
    input clk,
    input hidden_go,
    input reset,
    input signed [WIDTH*averaged_pixels_nr-1:0] hidden_in,
    output signed [4*WIDTH*HL_neurons-1:0] hidden_out,
    output hidden_done
    );
    
    wire signed [4*WIDTH*HL_neurons-1:0] dense_out;
    wire dense_done;
    
    //Biases and weights
    localparam signed [WIDTH*HL_neurons-1:0] biases_HL_param = { 8'sb11110111, 8'sb11110010, 8'sb00000001, 8'sb00000111, 8'sb00000100, 8'sb11111111, 8'sb00010011, 8'sb00001101, 8'sb11110100, 8'sb00010111, 8'sb00001010, 8'sb11111111, 8'sb11101011, 8'sb11111100, 8'sb00011111, 8'sb00010101, 8'sb11111011, 8'sb00001011, 8'sb00000011, 8'sb00001001, 8'sb00011100, 8'sb00010001, 8'sb00100100, 8'sb00001011, 8'sb00000011, 8'sb11111111, 8'sb11111111, 8'sb00100010, 8'sb00011000, 8'sb11111110, 8'sb00001101, 8'sb00001010 };
    
    localparam signed [WIDTH*HL_neurons*averaged_pixels_nr-1:0] weights_HL_param =   {
    8'sb11111100, 8'sb00001001, 8'sb00000111, 8'sb11111101, 8'sb00001010, 8'sb00001000, 8'sb00000010, 8'sb00000110, 8'sb00001011, 8'sb00000101, 8'sb11111101, 8'sb00001011, 8'sb00000011, 8'sb11111101, 8'sb11111001, 8'sb00000111, 8'sb00000010, 8'sb00001101, 8'sb00000100, 8'sb00000010, 8'sb11101110, 8'sb11100011, 8'sb11010000, 8'sb11010111, 8'sb11000010, 8'sb11111011, 8'sb11110100, 8'sb11111100, 8'sb11111111, 8'sb11100111, 8'sb11111110, 8'sb11111101, 8'sb00001000, 8'sb11111101, 8'sb11110111, 8'sb11110011, 8'sb11111101, 8'sb11110000, 8'sb11110100, 8'sb00001001, 8'sb11111110, 8'sb11111100, 8'sb00010101, 8'sb00000100, 8'sb00011110, 8'sb00001101, 8'sb00001011, 8'sb00010100, 8'sb00000001, 8'sb00000011, 8'sb00001011, 8'sb00001110, 8'sb00001110, 8'sb00011100, 8'sb00000010, 8'sb11100111, 8'sb00111001, 8'sb00011011, 8'sb00010101, 8'sb00010000, 8'sb00010010, 8'sb00010100, 8'sb00100010, 8'sb00101010, 8'sb00010011, 8'sb00010001, 8'sb00010101, 8'sb00100110, 8'sb11101110, 8'sb00001001, 8'sb00111110, 8'sb00000100, 8'sb00001110, 8'sb00010110, 8'sb00010001, 8'sb00100100, 8'sb11110010, 8'sb11100101, 8'sb00000101, 8'sb00000000, 8'sb11111111, 8'sb11110011, 8'sb11101000, 8'sb00100111, 8'sb00101001, 8'sb11111100, 8'sb00010100, 8'sb00011010, 8'sb00001011, 8'sb11000110, 8'sb10001000, 8'sb11010101, 8'sb11110111, 8'sb11111000, 8'sb11101010, 8'sb11100110, 8'sb11110111, 8'sb00110000, 8'sb00011001, 8'sb11101000, 8'sb11011111, 8'sb11010111, 8'sb10101011, 8'sb10111010, 8'sb11110000, 8'sb11100000, 8'sb11100000, 8'sb11100110, 8'sb11101001, 8'sb11011011, 8'sb11001111, 8'sb00100101, 8'sb11111101, 8'sb11100011, 8'sb11000111, 8'sb10100101, 8'sb10111001, 8'sb00001001, 8'sb00010101, 8'sb11110000, 8'sb11011110, 8'sb11011101, 8'sb11001110, 8'sb11100001, 8'sb11110110, 8'sb00110000, 8'sb00010011, 8'sb11100110, 8'sb11101011, 8'sb11101101, 8'sb00001000, 8'sb00011111, 8'sb00101100, 8'sb00000101, 8'sb11110001, 8'sb11101110, 8'sb11110110, 8'sb11111110, 8'sb00011000, 8'sb01000000, 8'sb00011100, 8'sb00011000, 8'sb00000000, 8'sb00000110, 8'sb00000001, 8'sb00011000, 8'sb00100011, 8'sb00101010, 8'sb00100101, 8'sb00011111, 8'sb00010010, 8'sb00010000, 8'sb00010010, 8'sb00110010, 8'sb11110010, 8'sb00000100, 8'sb00000100, 8'sb00000110, 8'sb00001101, 8'sb00001111, 8'sb00011001, 8'sb00100000, 8'sb00011100, 8'sb00101111, 8'sb00011111, 8'sb00101101, 8'sb00110010, 8'sb00011001, 8'sb11111000, 8'sb11100001, 8'sb11111101, 8'sb00001110, 8'sb00000001, 8'sb11111010, 8'sb00010111, 8'sb00011101, 8'sb00001111, 8'sb00100110, 8'sb00001001, 8'sb00011010, 8'sb00111100, 8'sb00010100, 8'sb11111000, 8'sb00001010, 8'sb11100000, 8'sb00011001, 8'sb00111101, 8'sb00000110, 8'sb00000000, 8'sb00010010, 8'sb11111001, 8'sb00011100, 8'sb11110110, 8'sb11110100, 8'sb00000110, 8'sb00000110,
    8'sb11111011, 8'sb00001001, 8'sb11111110, 8'sb00100011, 8'sb00110101, 8'sb00110011, 8'sb00101111, 8'sb11101000, 8'sb00111010, 8'sb01000001, 8'sb00101110, 8'sb00001110, 8'sb00000101, 8'sb00000101, 8'sb11111101, 8'sb00011001, 8'sb00000001, 8'sb00001101, 8'sb00101000, 8'sb00100110, 8'sb00010111, 8'sb00010001, 8'sb00000001, 8'sb11110000, 8'sb11111110, 8'sb00100101, 8'sb00001011, 8'sb00001100, 8'sb11111100, 8'sb11011100, 8'sb00000101, 8'sb00001100, 8'sb00000000, 8'sb00000011, 8'sb00010100, 8'sb00000110, 8'sb00010001, 8'sb11111010, 8'sb11111100, 8'sb11101010, 8'sb11100011, 8'sb00000101, 8'sb11010100, 8'sb11101110, 8'sb11101110, 8'sb11110000, 8'sb11110001, 8'sb00000010, 8'sb00000011, 8'sb00011000, 8'sb00011010, 8'sb11111010, 8'sb11111010, 8'sb00000011, 8'sb11111000, 8'sb11101100, 8'sb11111001, 8'sb11110110, 8'sb00000000, 8'sb11110011, 8'sb11111101, 8'sb00000100, 8'sb11110100, 8'sb11110110, 8'sb00000001, 8'sb00011010, 8'sb00001010, 8'sb00010111, 8'sb11111111, 8'sb11100011, 8'sb11110001, 8'sb11100111, 8'sb00010101, 8'sb00000110, 8'sb11111101, 8'sb11110110, 8'sb11111010, 8'sb11011000, 8'sb11100100, 8'sb00011010, 8'sb00100111, 8'sb00101000, 8'sb11111110, 8'sb11001111, 8'sb11110101, 8'sb00000010, 8'sb00011100, 8'sb00011111, 8'sb00000110, 8'sb11111001, 8'sb11100101, 8'sb11100101, 8'sb11101011, 8'sb00001111, 8'sb00011111, 8'sb01000100, 8'sb01001011, 8'sb11011011, 8'sb11100110, 8'sb11010100, 8'sb11111011, 8'sb00101101, 8'sb00100000, 8'sb00010100, 8'sb00001011, 8'sb00001000, 8'sb00001010, 8'sb00110010, 8'sb00110011, 8'sb00100100, 8'sb00100011, 8'sb00110011, 8'sb11101010, 8'sb11001010, 8'sb00000110, 8'sb00101100, 8'sb01000001, 8'sb00111000, 8'sb00010001, 8'sb00011000, 8'sb00010110, 8'sb00001110, 8'sb00010010, 8'sb00001010, 8'sb00010001, 8'sb00011110, 8'sb11111101, 8'sb11010000, 8'sb11110000, 8'sb00010010, 8'sb00011101, 8'sb00100111, 8'sb00001000, 8'sb00010111, 8'sb00001100, 8'sb11111110, 8'sb00000010, 8'sb11110111, 8'sb11101110, 8'sb00001101, 8'sb00010011, 8'sb00000110, 8'sb11111001, 8'sb11111011, 8'sb00001101, 8'sb00001011, 8'sb00000110, 8'sb00000110, 8'sb11110010, 8'sb11110011, 8'sb11101010, 8'sb11101100, 8'sb11100110, 8'sb00010001, 8'sb11110001, 8'sb00000100, 8'sb11100111, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00001010, 8'sb11110111, 8'sb11101000, 8'sb11011110, 8'sb11110100, 8'sb00001011, 8'sb11111011, 8'sb11010000, 8'sb00000011, 8'sb11010100, 8'sb11111110, 8'sb11111011, 8'sb11110111, 8'sb11111111, 8'sb11101010, 8'sb11110000, 8'sb11001000, 8'sb11100100, 8'sb11110010, 8'sb00000001, 8'sb11111111, 8'sb11111100, 8'sb11111101, 8'sb00010011, 8'sb00111101, 8'sb00111100, 8'sb00111000, 8'sb00010101, 8'sb00001011, 8'sb00011101, 8'sb11010100, 8'sb00000001, 8'sb00011010, 8'sb11111101, 8'sb00011001, 8'sb00000011,
    8'sb00001011, 8'sb00000111, 8'sb00000110, 8'sb11110101, 8'sb00000101, 8'sb11110110, 8'sb00001000, 8'sb11011000, 8'sb11010101, 8'sb11110010, 8'sb11100101, 8'sb11110010, 8'sb11110100, 8'sb11111010, 8'sb00001011, 8'sb11111010, 8'sb00011011, 8'sb11111011, 8'sb11110101, 8'sb11110111, 8'sb11111001, 8'sb11110111, 8'sb00010010, 8'sb00110101, 8'sb00110100, 8'sb00110001, 8'sb00000000, 8'sb00011100, 8'sb00000100, 8'sb11110000, 8'sb11101011, 8'sb11110110, 8'sb11101011, 8'sb11110000, 8'sb11111000, 8'sb11111101, 8'sb00010111, 8'sb00011001, 8'sb00011100, 8'sb00100110, 8'sb00110011, 8'sb00010100, 8'sb00001011, 8'sb11101111, 8'sb11110111, 8'sb11111101, 8'sb00000011, 8'sb00000001, 8'sb11111110, 8'sb00011000, 8'sb00011011, 8'sb00100100, 8'sb00010000, 8'sb00001001, 8'sb00110110, 8'sb00011000, 8'sb11011110, 8'sb11101001, 8'sb11010011, 8'sb11111101, 8'sb00000011, 8'sb00001001, 8'sb00001100, 8'sb11101101, 8'sb00000001, 8'sb00001111, 8'sb00011011, 8'sb00001010, 8'sb00111000, 8'sb00101000, 8'sb11011111, 8'sb11101001, 8'sb11101001, 8'sb11110100, 8'sb11111101, 8'sb00001001, 8'sb00010111, 8'sb11111100, 8'sb00000101, 8'sb11111110, 8'sb11110000, 8'sb11101010, 8'sb00111011, 8'sb00111010, 8'sb00000101, 8'sb11111000, 8'sb00000010, 8'sb11110000, 8'sb11101011, 8'sb00011001, 8'sb00010101, 8'sb00010100, 8'sb00010100, 8'sb00001101, 8'sb11110001, 8'sb11010100, 8'sb10111101, 8'sb11101011, 8'sb00011110, 8'sb11110100, 8'sb11111010, 8'sb11101010, 8'sb11110001, 8'sb00010011, 8'sb11111111, 8'sb00000100, 8'sb00011001, 8'sb00011000, 8'sb00000010, 8'sb11110101, 8'sb11010100, 8'sb10110111, 8'sb00000001, 8'sb11101100, 8'sb11111000, 8'sb00000110, 8'sb11101001, 8'sb11110000, 8'sb11110100, 8'sb11111101, 8'sb00010101, 8'sb00010010, 8'sb00000111, 8'sb11100101, 8'sb11010001, 8'sb10111010, 8'sb11110100, 8'sb00010000, 8'sb00001111, 8'sb00010110, 8'sb00000110, 8'sb00001101, 8'sb00000001, 8'sb00001001, 8'sb00000110, 8'sb11110000, 8'sb11100111, 8'sb11011001, 8'sb11011000, 8'sb11011001, 8'sb00001101, 8'sb11011101, 8'sb11111100, 8'sb11111001, 8'sb00000000, 8'sb00000100, 8'sb00001001, 8'sb00010000, 8'sb11111111, 8'sb11011010, 8'sb11010110, 8'sb11011101, 8'sb11101010, 8'sb11100001, 8'sb11111100, 8'sb00000101, 8'sb11101001, 8'sb11101101, 8'sb00000001, 8'sb00010011, 8'sb00011101, 8'sb00010100, 8'sb11110111, 8'sb11011110, 8'sb11010000, 8'sb11101001, 8'sb00000010, 8'sb00001110, 8'sb00000010, 8'sb01000000, 8'sb01001000, 8'sb00011010, 8'sb00101010, 8'sb00110110, 8'sb00110010, 8'sb00101001, 8'sb00001001, 8'sb11111100, 8'sb11111001, 8'sb00001000, 8'sb11110010, 8'sb11101001, 8'sb11111110, 8'sb11111010, 8'sb00011010, 8'sb11111000, 8'sb11110101, 8'sb00101001, 8'sb00100011, 8'sb11110110, 8'sb11111011, 8'sb11110001, 8'sb00000010, 8'sb00010110, 8'sb11111111, 8'sb00000010,
    8'sb11111001, 8'sb00000100, 8'sb11111111, 8'sb11101100, 8'sb11100001, 8'sb11001100, 8'sb11000011, 8'sb00000010, 8'sb00100000, 8'sb11011000, 8'sb11011000, 8'sb11101001, 8'sb11111000, 8'sb00001000, 8'sb00000101, 8'sb00001011, 8'sb11100011, 8'sb11111010, 8'sb11010001, 8'sb11100001, 8'sb00001011, 8'sb00011100, 8'sb00100100, 8'sb00011011, 8'sb00100101, 8'sb00001001, 8'sb11010111, 8'sb11110101, 8'sb00000000, 8'sb11101000, 8'sb11110100, 8'sb00011101, 8'sb00100010, 8'sb00101001, 8'sb00001001, 8'sb00000110, 8'sb00011100, 8'sb11111110, 8'sb00010100, 8'sb00010100, 8'sb11110111, 8'sb11110010, 8'sb11100101, 8'sb11011101, 8'sb00001000, 8'sb00011000, 8'sb00011110, 8'sb00000010, 8'sb11011001, 8'sb10111110, 8'sb11111110, 8'sb00000100, 8'sb11110110, 8'sb00001000, 8'sb00000011, 8'sb00001000, 8'sb11100100, 8'sb11111110, 8'sb00001100, 8'sb00001000, 8'sb00010010, 8'sb11111110, 8'sb11011110, 8'sb11010110, 8'sb00100011, 8'sb00001001, 8'sb00001111, 8'sb00000010, 8'sb00011000, 8'sb00001011, 8'sb11110010, 8'sb11110010, 8'sb00000110, 8'sb11110111, 8'sb00011011, 8'sb00001110, 8'sb11001010, 8'sb11010011, 8'sb00000111, 8'sb11111011, 8'sb11110111, 8'sb11100111, 8'sb11101000, 8'sb00010011, 8'sb00000110, 8'sb11110111, 8'sb00000101, 8'sb11111110, 8'sb11110110, 8'sb00011101, 8'sb00010011, 8'sb11101010, 8'sb11101111, 8'sb00001001, 8'sb00001101, 8'sb11110100, 8'sb11100000, 8'sb11101000, 8'sb11110000, 8'sb11111110, 8'sb00010110, 8'sb00011000, 8'sb00001000, 8'sb11111000, 8'sb00011011, 8'sb00010101, 8'sb00001100, 8'sb00000011, 8'sb11110000, 8'sb11111000, 8'sb11010000, 8'sb00001001, 8'sb11110001, 8'sb00010110, 8'sb00010101, 8'sb00000100, 8'sb11110110, 8'sb11101101, 8'sb00010001, 8'sb00001001, 8'sb11111000, 8'sb11100110, 8'sb11101010, 8'sb11011001, 8'sb11000111, 8'sb00011001, 8'sb11101111, 8'sb00010110, 8'sb00001101, 8'sb11111111, 8'sb11100111, 8'sb11111001, 8'sb00100111, 8'sb11111111, 8'sb11101001, 8'sb11101100, 8'sb11110100, 8'sb11110110, 8'sb11111101, 8'sb00101101, 8'sb11101110, 8'sb11111100, 8'sb11101111, 8'sb11100100, 8'sb11010101, 8'sb00011001, 8'sb00000111, 8'sb11111101, 8'sb00001101, 8'sb00000110, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00010100, 8'sb11111111, 8'sb00001110, 8'sb11101000, 8'sb11001111, 8'sb11011010, 8'sb11110010, 8'sb00001010, 8'sb00010111, 8'sb00010110, 8'sb00010001, 8'sb00100010, 8'sb00100010, 8'sb00001011, 8'sb00010000, 8'sb00000000, 8'sb00001111, 8'sb11101000, 8'sb11010101, 8'sb11010101, 8'sb11101100, 8'sb00001011, 8'sb00101010, 8'sb00100001, 8'sb00001111, 8'sb11110010, 8'sb11111110, 8'sb00001001, 8'sb00000100, 8'sb00000110, 8'sb11110111, 8'sb11100010, 8'sb11100100, 8'sb11010101, 8'sb11010010, 8'sb11010010, 8'sb11000110, 8'sb11010100, 8'sb11100110, 8'sb11100000, 8'sb11110010, 8'sb11111010, 8'sb00000110,
    8'sb11111010, 8'sb00000001, 8'sb00001010, 8'sb00010001, 8'sb00000101, 8'sb00001000, 8'sb00001101, 8'sb00011001, 8'sb00110101, 8'sb00011011, 8'sb00101101, 8'sb00001110, 8'sb11111100, 8'sb11111010, 8'sb00001100, 8'sb00001001, 8'sb00001010, 8'sb00100110, 8'sb00111100, 8'sb01001101, 8'sb00110101, 8'sb00100010, 8'sb00000110, 8'sb11110100, 8'sb11100011, 8'sb11110111, 8'sb00010000, 8'sb11101101, 8'sb11111000, 8'sb11111110, 8'sb00101011, 8'sb00010101, 8'sb00010110, 8'sb11110110, 8'sb11111001, 8'sb00000010, 8'sb00010001, 8'sb00001011, 8'sb00000000, 8'sb11111011, 8'sb11110111, 8'sb00000101, 8'sb00011001, 8'sb11111111, 8'sb00010000, 8'sb11110010, 8'sb11011101, 8'sb11100100, 8'sb11010000, 8'sb00001000, 8'sb00001110, 8'sb11110000, 8'sb11101011, 8'sb11111101, 8'sb00001110, 8'sb11110111, 8'sb00100100, 8'sb00100100, 8'sb00100000, 8'sb11111110, 8'sb11111010, 8'sb11110010, 8'sb11100110, 8'sb00001001, 8'sb00010100, 8'sb11110101, 8'sb11111101, 8'sb11110001, 8'sb11010011, 8'sb11110100, 8'sb00100110, 8'sb00010011, 8'sb00001010, 8'sb00001010, 8'sb00001011, 8'sb11011111, 8'sb11011001, 8'sb00100000, 8'sb00000101, 8'sb11110110, 8'sb00001011, 8'sb00000000, 8'sb11101010, 8'sb11011110, 8'sb11101101, 8'sb11011110, 8'sb11101001, 8'sb11100101, 8'sb11100101, 8'sb11101001, 8'sb00101010, 8'sb00011101, 8'sb11110000, 8'sb11100011, 8'sb00000000, 8'sb11111000, 8'sb01011000, 8'sb00100110, 8'sb11101101, 8'sb11111111, 8'sb11101100, 8'sb11100101, 8'sb11110110, 8'sb00000110, 8'sb00111100, 8'sb00101100, 8'sb11110010, 8'sb11101100, 8'sb11100010, 8'sb00000000, 8'sb00110011, 8'sb01000001, 8'sb00001011, 8'sb00101101, 8'sb11111101, 8'sb00001110, 8'sb00011101, 8'sb00101010, 8'sb00100010, 8'sb00010011, 8'sb00001011, 8'sb00000110, 8'sb11110110, 8'sb00010100, 8'sb00111001, 8'sb00110010, 8'sb11101011, 8'sb00001101, 8'sb00001011, 8'sb00010001, 8'sb00100010, 8'sb00001010, 8'sb11111010, 8'sb00001010, 8'sb00011110, 8'sb00011001, 8'sb00010101, 8'sb00101011, 8'sb00100100, 8'sb00111001, 8'sb11101101, 8'sb00100000, 8'sb00001100, 8'sb00010111, 8'sb00001110, 8'sb11101100, 8'sb11110101, 8'sb00000111, 8'sb00011010, 8'sb00010111, 8'sb00011110, 8'sb11111110, 8'sb11011100, 8'sb00100011, 8'sb00001111, 8'sb00110101, 8'sb00011100, 8'sb00001010, 8'sb00000001, 8'sb00000011, 8'sb11111000, 8'sb11111101, 8'sb11110111, 8'sb11111110, 8'sb00000101, 8'sb11011011, 8'sb11001010, 8'sb11110001, 8'sb00000001, 8'sb11011001, 8'sb11011111, 8'sb11101001, 8'sb11111110, 8'sb11111101, 8'sb11101011, 8'sb11100010, 8'sb11100000, 8'sb11100101, 8'sb11101100, 8'sb11001101, 8'sb11111111, 8'sb00001000, 8'sb11111011, 8'sb11110011, 8'sb11011010, 8'sb11011010, 8'sb11000110, 8'sb11000010, 8'sb10011101, 8'sb10001011, 8'sb10011100, 8'sb11001010, 8'sb10100011, 8'sb11001110, 8'sb11110011, 8'sb11111001,
    8'sb11110110, 8'sb11110110, 8'sb00000111, 8'sb00100101, 8'sb00100000, 8'sb01000001, 8'sb00110001, 8'sb00000100, 8'sb00011110, 8'sb00111010, 8'sb00110100, 8'sb00010001, 8'sb00000110, 8'sb11110110, 8'sb00000010, 8'sb00001111, 8'sb00100101, 8'sb00001100, 8'sb11110110, 8'sb00001101, 8'sb00000111, 8'sb00101001, 8'sb00010111, 8'sb00011100, 8'sb00010100, 8'sb00100010, 8'sb11110110, 8'sb00000010, 8'sb00001011, 8'sb11001100, 8'sb11011110, 8'sb11110011, 8'sb00010011, 8'sb11110001, 8'sb11110011, 8'sb00000010, 8'sb00000010, 8'sb00001110, 8'sb00000101, 8'sb11110000, 8'sb11110001, 8'sb00011010, 8'sb11110001, 8'sb11001111, 8'sb11011100, 8'sb11111001, 8'sb00000101, 8'sb00000010, 8'sb11111010, 8'sb11110100, 8'sb11110011, 8'sb11101011, 8'sb00000110, 8'sb00001010, 8'sb00000100, 8'sb11110111, 8'sb11100110, 8'sb11100011, 8'sb11110101, 8'sb11111011, 8'sb00010100, 8'sb00000101, 8'sb11100110, 8'sb11101010, 8'sb11100110, 8'sb11111011, 8'sb00000111, 8'sb11101101, 8'sb11100010, 8'sb11101110, 8'sb11101111, 8'sb11001010, 8'sb11010111, 8'sb00001010, 8'sb00011001, 8'sb00001000, 8'sb11100011, 8'sb11011010, 8'sb11101100, 8'sb11111001, 8'sb00001101, 8'sb00001000, 8'sb11010101, 8'sb10111100, 8'sb11110011, 8'sb11000000, 8'sb11011011, 8'sb00001111, 8'sb00010111, 8'sb00011101, 8'sb11110011, 8'sb11110111, 8'sb00001101, 8'sb00001101, 8'sb00010111, 8'sb00100000, 8'sb11101111, 8'sb10101110, 8'sb00000001, 8'sb11011001, 8'sb11101000, 8'sb11111011, 8'sb11111110, 8'sb00010010, 8'sb00001111, 8'sb00001010, 8'sb00010000, 8'sb00000100, 8'sb11101101, 8'sb00000011, 8'sb11101100, 8'sb11010000, 8'sb11100111, 8'sb11010111, 8'sb10111111, 8'sb11010000, 8'sb11100100, 8'sb00010110, 8'sb00011000, 8'sb00010101, 8'sb00010101, 8'sb11110101, 8'sb11110001, 8'sb11110011, 8'sb00000111, 8'sb11000011, 8'sb11011111, 8'sb11010001, 8'sb10110101, 8'sb10101100, 8'sb11101010, 8'sb00110011, 8'sb00101111, 8'sb00000011, 8'sb00000000, 8'sb00000100, 8'sb11101010, 8'sb11111110, 8'sb11111100, 8'sb11010111, 8'sb00001111, 8'sb11001011, 8'sb10111011, 8'sb10101110, 8'sb11100011, 8'sb00011011, 8'sb00011101, 8'sb00100001, 8'sb00010010, 8'sb00000000, 8'sb11110010, 8'sb11111111, 8'sb11101110, 8'sb00000110, 8'sb11101100, 8'sb11101101, 8'sb11011001, 8'sb11010000, 8'sb11100000, 8'sb11100011, 8'sb00001101, 8'sb00010111, 8'sb00010101, 8'sb00001011, 8'sb00000101, 8'sb11111000, 8'sb11100000, 8'sb11110001, 8'sb00000100, 8'sb11011100, 8'sb11101011, 8'sb11010011, 8'sb11010010, 8'sb11110010, 8'sb11100111, 8'sb00000111, 8'sb00000010, 8'sb00001000, 8'sb11111110, 8'sb00000100, 8'sb11101101, 8'sb11100100, 8'sb11111001, 8'sb00001011, 8'sb00010000, 8'sb00011100, 8'sb00001110, 8'sb11111010, 8'sb00000110, 8'sb11110100, 8'sb11111011, 8'sb11111111, 8'sb11100101, 8'sb11100011, 8'sb11111111, 8'sb11111111,
    8'sb11111111, 8'sb11110101, 8'sb00001110, 8'sb00000111, 8'sb00011001, 8'sb00011111, 8'sb00100000, 8'sb11111111, 8'sb11011111, 8'sb00110000, 8'sb00110100, 8'sb00001111, 8'sb00000101, 8'sb00001000, 8'sb00001000, 8'sb00011111, 8'sb00001011, 8'sb00011100, 8'sb11101101, 8'sb11101110, 8'sb11010010, 8'sb11010010, 8'sb11110001, 8'sb00001100, 8'sb00011110, 8'sb00010101, 8'sb11110101, 8'sb00000011, 8'sb00000000, 8'sb00000101, 8'sb00001110, 8'sb11101011, 8'sb11101101, 8'sb11100101, 8'sb11010000, 8'sb11010110, 8'sb11011111, 8'sb11100111, 8'sb11101001, 8'sb00010111, 8'sb11110010, 8'sb11100111, 8'sb11001110, 8'sb11101011, 8'sb00000101, 8'sb11011100, 8'sb11110101, 8'sb11100100, 8'sb11100101, 8'sb11111110, 8'sb00000011, 8'sb11111001, 8'sb11111101, 8'sb00100001, 8'sb00001010, 8'sb00000001, 8'sb11010101, 8'sb11010011, 8'sb11100100, 8'sb11011101, 8'sb11101101, 8'sb11011110, 8'sb11111101, 8'sb00000100, 8'sb00001011, 8'sb11101011, 8'sb11110100, 8'sb11100110, 8'sb11100001, 8'sb11011010, 8'sb00010000, 8'sb11001111, 8'sb11000000, 8'sb11010111, 8'sb11110011, 8'sb11110101, 8'sb00011010, 8'sb00001101, 8'sb00000100, 8'sb11100000, 8'sb11011111, 8'sb11100010, 8'sb11000000, 8'sb11001110, 8'sb11110111, 8'sb11010101, 8'sb10100111, 8'sb11110101, 8'sb00001101, 8'sb00101001, 8'sb01000100, 8'sb00100000, 8'sb00010000, 8'sb00001011, 8'sb11111101, 8'sb11101000, 8'sb11000000, 8'sb11000000, 8'sb11111011, 8'sb00000000, 8'sb11010010, 8'sb11010010, 8'sb00011001, 8'sb00111010, 8'sb00101001, 8'sb00001101, 8'sb00011111, 8'sb00001110, 8'sb11111010, 8'sb11001010, 8'sb10111100, 8'sb10111110, 8'sb00010000, 8'sb11011110, 8'sb11011000, 8'sb11010000, 8'sb00000011, 8'sb00100001, 8'sb00001001, 8'sb11111101, 8'sb00000001, 8'sb00000000, 8'sb11110100, 8'sb11011001, 8'sb11000001, 8'sb11001100, 8'sb11110010, 8'sb11011001, 8'sb11001111, 8'sb11011110, 8'sb11101111, 8'sb00000001, 8'sb00010110, 8'sb00000101, 8'sb11111100, 8'sb11110001, 8'sb11010011, 8'sb11011011, 8'sb11011111, 8'sb11110111, 8'sb00001110, 8'sb11110010, 8'sb11101001, 8'sb11100001, 8'sb11011110, 8'sb11101110, 8'sb11111101, 8'sb00000011, 8'sb11111000, 8'sb11101011, 8'sb11010100, 8'sb11101000, 8'sb11101001, 8'sb00001100, 8'sb00010101, 8'sb11011100, 8'sb00001011, 8'sb11111100, 8'sb00000111, 8'sb11110110, 8'sb11101100, 8'sb11101100, 8'sb11110101, 8'sb00001101, 8'sb11110000, 8'sb11110101, 8'sb11111001, 8'sb00100010, 8'sb11111101, 8'sb11100001, 8'sb00001101, 8'sb11111111, 8'sb00001001, 8'sb11110100, 8'sb11101101, 8'sb11111001, 8'sb00000101, 8'sb00010111, 8'sb00000000, 8'sb00100010, 8'sb00001011, 8'sb11111010, 8'sb11111110, 8'sb00010001, 8'sb00010110, 8'sb00001100, 8'sb11111110, 8'sb00000000, 8'sb11101100, 8'sb00010010, 8'sb00010000, 8'sb11011011, 8'sb11101111, 8'sb11011110, 8'sb00000101, 8'sb00000001,
    8'sb11111110, 8'sb00001011, 8'sb11111010, 8'sb11101110, 8'sb11110010, 8'sb11010101, 8'sb11011101, 8'sb11100001, 8'sb11010011, 8'sb11100110, 8'sb11101000, 8'sb11101100, 8'sb00000000, 8'sb00000111, 8'sb00001100, 8'sb00000011, 8'sb11111101, 8'sb11011100, 8'sb11000011, 8'sb10110100, 8'sb10111101, 8'sb10111000, 8'sb11000111, 8'sb11010001, 8'sb11001010, 8'sb11110110, 8'sb00010000, 8'sb00000000, 8'sb11111111, 8'sb11011111, 8'sb00100001, 8'sb00010001, 8'sb00001010, 8'sb11110000, 8'sb11110111, 8'sb11110001, 8'sb11101011, 8'sb11110011, 8'sb11110111, 8'sb00000000, 8'sb11111110, 8'sb00001101, 8'sb11101010, 8'sb00010000, 8'sb11111101, 8'sb00011111, 8'sb00010011, 8'sb11111011, 8'sb11101111, 8'sb11111000, 8'sb00001000, 8'sb11101101, 8'sb00001001, 8'sb11111110, 8'sb11101000, 8'sb11111000, 8'sb00100000, 8'sb00010010, 8'sb00010110, 8'sb00010100, 8'sb00000001, 8'sb00001100, 8'sb00000101, 8'sb00010001, 8'sb00000101, 8'sb00000110, 8'sb11100011, 8'sb11010110, 8'sb11101010, 8'sb00001101, 8'sb00111000, 8'sb00000101, 8'sb00010111, 8'sb00001101, 8'sb00010010, 8'sb00011000, 8'sb00001110, 8'sb00101011, 8'sb00101100, 8'sb00000111, 8'sb11001111, 8'sb11010101, 8'sb11010110, 8'sb11101100, 8'sb00111101, 8'sb00110100, 8'sb11111100, 8'sb00000000, 8'sb00010001, 8'sb00010010, 8'sb11110101, 8'sb00100011, 8'sb00101100, 8'sb00001110, 8'sb11101000, 8'sb11110110, 8'sb11010010, 8'sb11001100, 8'sb00000011, 8'sb00011110, 8'sb00000011, 8'sb11100010, 8'sb11101000, 8'sb11101111, 8'sb11111111, 8'sb00100011, 8'sb00100101, 8'sb00000010, 8'sb11011101, 8'sb11110100, 8'sb11100001, 8'sb11001111, 8'sb00001000, 8'sb11100101, 8'sb11000001, 8'sb11000111, 8'sb11001100, 8'sb11101111, 8'sb00010100, 8'sb00101100, 8'sb00001111, 8'sb11010110, 8'sb11100000, 8'sb11011111, 8'sb11110000, 8'sb11110011, 8'sb00100000, 8'sb11101101, 8'sb10100010, 8'sb10000001, 8'sb11010111, 8'sb00010001, 8'sb00101101, 8'sb00001000, 8'sb11010110, 8'sb11100011, 8'sb11101101, 8'sb10111111, 8'sb11110110, 8'sb00100100, 8'sb00001000, 8'sb11000100, 8'sb10010111, 8'sb10101111, 8'sb11101010, 8'sb00000110, 8'sb00000111, 8'sb00000100, 8'sb11111110, 8'sb11111001, 8'sb11101111, 8'sb11011011, 8'sb11110010, 8'sb00000001, 8'sb00000110, 8'sb11000110, 8'sb11001110, 8'sb11100001, 8'sb11110000, 8'sb11110100, 8'sb00001000, 8'sb00001110, 8'sb00001101, 8'sb00000110, 8'sb00000111, 8'sb11101110, 8'sb00001110, 8'sb00010000, 8'sb11111100, 8'sb11100011, 8'sb11100110, 8'sb11110000, 8'sb11001100, 8'sb11100110, 8'sb11101101, 8'sb00000010, 8'sb11110100, 8'sb00001001, 8'sb11111111, 8'sb11110010, 8'sb11101010, 8'sb00000010, 8'sb11110100, 8'sb00000010, 8'sb11110010, 8'sb00100001, 8'sb00101100, 8'sb11111110, 8'sb11110101, 8'sb11101011, 8'sb11111000, 8'sb00000000, 8'sb11110101, 8'sb11111111, 8'sb11111010, 8'sb11111011,
    8'sb00000010, 8'sb11111010, 8'sb00000010, 8'sb11110011, 8'sb11110001, 8'sb11011001, 8'sb11010001, 8'sb11011110, 8'sb00011000, 8'sb11010111, 8'sb11011101, 8'sb11101000, 8'sb11111000, 8'sb11111001, 8'sb00000101, 8'sb00000010, 8'sb11110110, 8'sb00001100, 8'sb00011000, 8'sb00001100, 8'sb11100101, 8'sb11001100, 8'sb11011001, 8'sb11110010, 8'sb11111110, 8'sb00000010, 8'sb00100000, 8'sb11111010, 8'sb11111100, 8'sb11110101, 8'sb11101110, 8'sb00000010, 8'sb00001001, 8'sb00100010, 8'sb00011110, 8'sb00001111, 8'sb11101111, 8'sb11101011, 8'sb11111001, 8'sb11101101, 8'sb00010000, 8'sb00010001, 8'sb11110010, 8'sb00100110, 8'sb11110000, 8'sb00000010, 8'sb00010100, 8'sb00011010, 8'sb00100110, 8'sb00101001, 8'sb00010101, 8'sb00000001, 8'sb11111001, 8'sb11011011, 8'sb11110001, 8'sb11110101, 8'sb00000011, 8'sb00010101, 8'sb00011000, 8'sb00011100, 8'sb00011000, 8'sb00000111, 8'sb00010010, 8'sb00011110, 8'sb00011111, 8'sb00001101, 8'sb11110011, 8'sb11110000, 8'sb11111001, 8'sb00101011, 8'sb00000001, 8'sb00001011, 8'sb00101101, 8'sb00100110, 8'sb00000100, 8'sb00010010, 8'sb00000101, 8'sb00011000, 8'sb00010010, 8'sb00011101, 8'sb00001100, 8'sb11101111, 8'sb00010100, 8'sb00110010, 8'sb00010110, 8'sb00000101, 8'sb00000100, 8'sb11011101, 8'sb11100010, 8'sb11010000, 8'sb11011100, 8'sb00000110, 8'sb00010111, 8'sb00101001, 8'sb11111001, 8'sb11110000, 8'sb11111011, 8'sb00010011, 8'sb11101101, 8'sb00000011, 8'sb10111011, 8'sb11000111, 8'sb11001010, 8'sb11110001, 8'sb11111010, 8'sb00001100, 8'sb00011001, 8'sb00000011, 8'sb11010010, 8'sb11011011, 8'sb11010111, 8'sb00001101, 8'sb00000101, 8'sb00000000, 8'sb10111011, 8'sb11011101, 8'sb00010010, 8'sb00001110, 8'sb00000011, 8'sb00000010, 8'sb00000111, 8'sb11100101, 8'sb11110101, 8'sb11111001, 8'sb11111011, 8'sb00010110, 8'sb00010101, 8'sb11100101, 8'sb10111101, 8'sb00000010, 8'sb00011010, 8'sb00011010, 8'sb00001000, 8'sb00001010, 8'sb11111101, 8'sb11110100, 8'sb11110110, 8'sb11111100, 8'sb00001100, 8'sb00100111, 8'sb11110111, 8'sb11111110, 8'sb11100101, 8'sb00000011, 8'sb00001001, 8'sb11111011, 8'sb11111100, 8'sb11110000, 8'sb11110010, 8'sb11100110, 8'sb11111100, 8'sb11111111, 8'sb00001011, 8'sb11100010, 8'sb11110001, 8'sb11101110, 8'sb11100010, 8'sb00000001, 8'sb00000100, 8'sb00000100, 8'sb00000010, 8'sb11110111, 8'sb11110011, 8'sb11111010, 8'sb00000011, 8'sb00011111, 8'sb00001010, 8'sb11011101, 8'sb00000010, 8'sb11011111, 8'sb00001110, 8'sb00010000, 8'sb00001001, 8'sb11111101, 8'sb00000111, 8'sb00010110, 8'sb00010010, 8'sb00011101, 8'sb00010001, 8'sb11111010, 8'sb11111101, 8'sb11111011, 8'sb00000111, 8'sb00011010, 8'sb00011010, 8'sb01000111, 8'sb01101001, 8'sb01001011, 8'sb01001000, 8'sb01001100, 8'sb01000000, 8'sb00111011, 8'sb01001101, 8'sb00110011, 8'sb11111001, 8'sb00000010,
    8'sb11111100, 8'sb11111000, 8'sb00000001, 8'sb00000011, 8'sb00001110, 8'sb00000011, 8'sb11110001, 8'sb00000101, 8'sb00100101, 8'sb11010110, 8'sb11100010, 8'sb11111100, 8'sb11111001, 8'sb00001000, 8'sb11111010, 8'sb00000111, 8'sb11111110, 8'sb11101110, 8'sb00001000, 8'sb11110110, 8'sb00000110, 8'sb11110101, 8'sb00001000, 8'sb11101100, 8'sb11001001, 8'sb11010010, 8'sb11011000, 8'sb00001110, 8'sb11110101, 8'sb11101000, 8'sb11011010, 8'sb11001101, 8'sb11011010, 8'sb11110001, 8'sb11101100, 8'sb11101000, 8'sb11010010, 8'sb10100000, 8'sb10110101, 8'sb11000000, 8'sb11010001, 8'sb11110110, 8'sb00010011, 8'sb11101001, 8'sb11100011, 8'sb11110110, 8'sb11010110, 8'sb11100011, 8'sb11100111, 8'sb11101101, 8'sb11101001, 8'sb11100100, 8'sb11101111, 8'sb00001000, 8'sb11111001, 8'sb00001011, 8'sb00110010, 8'sb00001010, 8'sb11011010, 8'sb11011111, 8'sb11011010, 8'sb11111000, 8'sb00000010, 8'sb00010111, 8'sb00111000, 8'sb00111011, 8'sb00110101, 8'sb00110100, 8'sb00110100, 8'sb00001111, 8'sb00010000, 8'sb00010100, 8'sb11000110, 8'sb11111100, 8'sb11111110, 8'sb00001011, 8'sb00011001, 8'sb00010011, 8'sb00001001, 8'sb00010010, 8'sb00100010, 8'sb00111011, 8'sb01001101, 8'sb01000000, 8'sb11111000, 8'sb11110011, 8'sb11101000, 8'sb11110100, 8'sb00010001, 8'sb00011101, 8'sb00011010, 8'sb11110111, 8'sb11011011, 8'sb11000110, 8'sb11000101, 8'sb11010101, 8'sb00001100, 8'sb01000111, 8'sb00000101, 8'sb11011001, 8'sb00000110, 8'sb00000000, 8'sb00010000, 8'sb00011011, 8'sb00000001, 8'sb11111100, 8'sb00000110, 8'sb11110100, 8'sb11010110, 8'sb11001101, 8'sb11111101, 8'sb00011101, 8'sb11110011, 8'sb11110010, 8'sb00011011, 8'sb00011100, 8'sb00010001, 8'sb00001111, 8'sb11111100, 8'sb00000011, 8'sb00001010, 8'sb11110100, 8'sb11100110, 8'sb11101001, 8'sb00000100, 8'sb00011100, 8'sb00101001, 8'sb11010000, 8'sb00000010, 8'sb00010110, 8'sb00100001, 8'sb00010010, 8'sb00000100, 8'sb11111111, 8'sb11111011, 8'sb00001011, 8'sb11110100, 8'sb00001101, 8'sb00000101, 8'sb11101100, 8'sb00001011, 8'sb11011001, 8'sb11111000, 8'sb11110001, 8'sb11110000, 8'sb11101101, 8'sb11101110, 8'sb11100111, 8'sb11110100, 8'sb11111110, 8'sb00011010, 8'sb00000001, 8'sb00101001, 8'sb11111110, 8'sb11111101, 8'sb00001011, 8'sb00001100, 8'sb11111100, 8'sb11111001, 8'sb11110111, 8'sb11111000, 8'sb11101110, 8'sb11101111, 8'sb11101010, 8'sb11111010, 8'sb00011110, 8'sb00111101, 8'sb00000110, 8'sb00000111, 8'sb00001101, 8'sb11101111, 8'sb10111100, 8'sb11100100, 8'sb11111111, 8'sb11100110, 8'sb11111000, 8'sb00000100, 8'sb00001000, 8'sb00001001, 8'sb00010100, 8'sb00100011, 8'sb11110101, 8'sb11110101, 8'sb11111110, 8'sb11101100, 8'sb11010001, 8'sb11001100, 8'sb11111101, 8'sb00000110, 8'sb11111100, 8'sb00010100, 8'sb00000110, 8'sb00001111, 8'sb00010101, 8'sb11111010, 8'sb00000011,
    8'sb00000001, 8'sb11111111, 8'sb11111010, 8'sb11101101, 8'sb11101010, 8'sb11110001, 8'sb11100010, 8'sb11111011, 8'sb11011101, 8'sb11100111, 8'sb11100011, 8'sb00000010, 8'sb00001010, 8'sb11111101, 8'sb00001000, 8'sb00000110, 8'sb11110001, 8'sb11001101, 8'sb11000111, 8'sb11000000, 8'sb10110101, 8'sb11010011, 8'sb11110101, 8'sb00010101, 8'sb11111000, 8'sb11110100, 8'sb11111010, 8'sb11111101, 8'sb00010111, 8'sb00011000, 8'sb00010011, 8'sb00001000, 8'sb11101111, 8'sb00000000, 8'sb00001010, 8'sb11111101, 8'sb00100001, 8'sb00011101, 8'sb00001001, 8'sb00000101, 8'sb00001100, 8'sb00000011, 8'sb00010010, 8'sb00000001, 8'sb00010101, 8'sb00001011, 8'sb00001101, 8'sb00000010, 8'sb00001011, 8'sb11111011, 8'sb00001000, 8'sb11101111, 8'sb11111100, 8'sb11111001, 8'sb11101110, 8'sb11111011, 8'sb11011001, 8'sb00100101, 8'sb00100110, 8'sb00011011, 8'sb00001010, 8'sb11110111, 8'sb11111110, 8'sb11110001, 8'sb00001111, 8'sb00010000, 8'sb00001010, 8'sb00001100, 8'sb11111001, 8'sb11110001, 8'sb11100110, 8'sb00101100, 8'sb11111000, 8'sb00000110, 8'sb11110000, 8'sb11101111, 8'sb11101110, 8'sb00000001, 8'sb00010100, 8'sb00001001, 8'sb11111110, 8'sb11111110, 8'sb11011110, 8'sb11100011, 8'sb11100100, 8'sb00000010, 8'sb11111100, 8'sb00010100, 8'sb00001001, 8'sb00100100, 8'sb00011111, 8'sb00011111, 8'sb00011011, 8'sb11110100, 8'sb11111111, 8'sb11111011, 8'sb11111000, 8'sb00000011, 8'sb00001110, 8'sb00001111, 8'sb11110000, 8'sb11111000, 8'sb00001110, 8'sb00010011, 8'sb00110001, 8'sb00111001, 8'sb00010101, 8'sb11110011, 8'sb00000011, 8'sb00001001, 8'sb11110001, 8'sb11111001, 8'sb00100011, 8'sb00000011, 8'sb11001011, 8'sb11010100, 8'sb11100011, 8'sb11010101, 8'sb00100000, 8'sb00101100, 8'sb00000101, 8'sb11100000, 8'sb11110100, 8'sb11111110, 8'sb00001001, 8'sb11011101, 8'sb11011110, 8'sb00000110, 8'sb11101001, 8'sb11100100, 8'sb10111100, 8'sb11000101, 8'sb11000001, 8'sb11100101, 8'sb11110011, 8'sb11110010, 8'sb11111000, 8'sb11111101, 8'sb11010011, 8'sb11111010, 8'sb00010010, 8'sb00010100, 8'sb00001010, 8'sb00000101, 8'sb11101100, 8'sb11100101, 8'sb11010100, 8'sb00000100, 8'sb11111111, 8'sb00000001, 8'sb00000110, 8'sb00001100, 8'sb11011011, 8'sb11110111, 8'sb11111101, 8'sb00110000, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00001010, 8'sb00001000, 8'sb00010001, 8'sb00001011, 8'sb00001001, 8'sb00001100, 8'sb11111111, 8'sb11011100, 8'sb00010110, 8'sb11110110, 8'sb00101000, 8'sb00101010, 8'sb00101100, 8'sb00100000, 8'sb00011011, 8'sb00000011, 8'sb00001000, 8'sb11101010, 8'sb11110001, 8'sb11111101, 8'sb11100111, 8'sb11000100, 8'sb11111110, 8'sb11111111, 8'sb11110100, 8'sb00001000, 8'sb00011001, 8'sb00101101, 8'sb00010000, 8'sb11111110, 8'sb11111001, 8'sb00000001, 8'sb11010000, 8'sb11001011, 8'sb11101010, 8'sb11110111, 8'sb11111010,
    8'sb00001001, 8'sb00001001, 8'sb11111001, 8'sb00000111, 8'sb11110000, 8'sb11101001, 8'sb11101011, 8'sb00010011, 8'sb00010010, 8'sb11101101, 8'sb11101000, 8'sb11110101, 8'sb00000010, 8'sb00000011, 8'sb00000100, 8'sb11101110, 8'sb11101111, 8'sb00000100, 8'sb00010001, 8'sb00100110, 8'sb00111100, 8'sb01000011, 8'sb00110010, 8'sb00000101, 8'sb11100001, 8'sb11100010, 8'sb11100001, 8'sb11101011, 8'sb11111101, 8'sb11110101, 8'sb00000000, 8'sb11110010, 8'sb00000101, 8'sb11110100, 8'sb11111101, 8'sb00100111, 8'sb00110011, 8'sb00101101, 8'sb00001010, 8'sb11110110, 8'sb10111100, 8'sb11001110, 8'sb00110010, 8'sb00100000, 8'sb11110011, 8'sb11101000, 8'sb11111100, 8'sb00000101, 8'sb00010011, 8'sb00010000, 8'sb00101100, 8'sb00101110, 8'sb00011001, 8'sb00000011, 8'sb11000101, 8'sb11011001, 8'sb00111110, 8'sb00010001, 8'sb11110110, 8'sb00001100, 8'sb00010001, 8'sb00000110, 8'sb11010011, 8'sb11010110, 8'sb00111001, 8'sb00110000, 8'sb00010110, 8'sb00001011, 8'sb10001101, 8'sb10111011, 8'sb00010011, 8'sb11101010, 8'sb11100010, 8'sb11011011, 8'sb11001110, 8'sb11010000, 8'sb10111000, 8'sb11000001, 8'sb00100111, 8'sb00100110, 8'sb00100011, 8'sb11111101, 8'sb10101011, 8'sb11010101, 8'sb00000111, 8'sb11011000, 8'sb11001110, 8'sb11100110, 8'sb11111010, 8'sb00000001, 8'sb11101100, 8'sb11100010, 8'sb11111100, 8'sb00001110, 8'sb11111110, 8'sb11100001, 8'sb11100010, 8'sb11110010, 8'sb00001110, 8'sb00001110, 8'sb00000110, 8'sb00100110, 8'sb00001010, 8'sb11111111, 8'sb11111000, 8'sb11110000, 8'sb00010000, 8'sb11110100, 8'sb11101100, 8'sb11100110, 8'sb11110000, 8'sb00001111, 8'sb00101001, 8'sb00010000, 8'sb00011001, 8'sb11111000, 8'sb11111001, 8'sb00000100, 8'sb11110011, 8'sb11101000, 8'sb11111011, 8'sb11101011, 8'sb11100000, 8'sb11110101, 8'sb11111001, 8'sb00100010, 8'sb00010101, 8'sb00001011, 8'sb00000100, 8'sb11111011, 8'sb00011100, 8'sb00001111, 8'sb00010001, 8'sb11111011, 8'sb00010000, 8'sb00001000, 8'sb11101010, 8'sb11111101, 8'sb11111101, 8'sb00110011, 8'sb00100010, 8'sb00100100, 8'sb00000101, 8'sb00001110, 8'sb00001011, 8'sb00010111, 8'sb00001010, 8'sb11110101, 8'sb11111010, 8'sb00000001, 8'sb00000110, 8'sb00000101, 8'sb00000010, 8'sb00100110, 8'sb00000110, 8'sb00001000, 8'sb00010001, 8'sb00010110, 8'sb00000100, 8'sb00001001, 8'sb00000000, 8'sb11111111, 8'sb11111100, 8'sb00000110, 8'sb11110101, 8'sb00000110, 8'sb00000010, 8'sb11111101, 8'sb00000000, 8'sb00011000, 8'sb00011101, 8'sb00000010, 8'sb00001010, 8'sb00011001, 8'sb00010110, 8'sb00000111, 8'sb11111101, 8'sb11100000, 8'sb11011111, 8'sb11100110, 8'sb11111000, 8'sb11111011, 8'sb00001000, 8'sb11101100, 8'sb11101001, 8'sb00000000, 8'sb00010100, 8'sb00001101, 8'sb11111110, 8'sb00100110, 8'sb00101101, 8'sb11101111, 8'sb11101000, 8'sb11111000, 8'sb11111000, 8'sb11111101,
    8'sb00000010, 8'sb00001010, 8'sb11111111, 8'sb00000101, 8'sb00011100, 8'sb00011101, 8'sb00010100, 8'sb00000110, 8'sb00011100, 8'sb00010011, 8'sb00001110, 8'sb00001111, 8'sb00000010, 8'sb00001010, 8'sb00000000, 8'sb00001010, 8'sb11101111, 8'sb11111101, 8'sb00101000, 8'sb00011100, 8'sb00000010, 8'sb11111100, 8'sb00000110, 8'sb00010000, 8'sb00010000, 8'sb00011100, 8'sb00100011, 8'sb00011010, 8'sb11111100, 8'sb11100111, 8'sb10111101, 8'sb11110001, 8'sb11100111, 8'sb00010101, 8'sb00011110, 8'sb00100011, 8'sb00101110, 8'sb00100111, 8'sb00001110, 8'sb11111100, 8'sb00001010, 8'sb00110010, 8'sb11101001, 8'sb11010001, 8'sb11100101, 8'sb11101111, 8'sb00001010, 8'sb00010011, 8'sb00011101, 8'sb00101011, 8'sb00011010, 8'sb11111111, 8'sb00001010, 8'sb00001011, 8'sb00001101, 8'sb11110010, 8'sb11110101, 8'sb11101011, 8'sb11111010, 8'sb00000010, 8'sb00010110, 8'sb00001100, 8'sb00000101, 8'sb11100011, 8'sb11110001, 8'sb00000000, 8'sb11111001, 8'sb11111101, 8'sb00010100, 8'sb00001110, 8'sb11011101, 8'sb11100101, 8'sb11110011, 8'sb00011010, 8'sb00010110, 8'sb11110111, 8'sb11100110, 8'sb11011010, 8'sb11111101, 8'sb00001000, 8'sb11110011, 8'sb11101110, 8'sb00011100, 8'sb00001101, 8'sb11100000, 8'sb00000011, 8'sb11110011, 8'sb11111111, 8'sb00000011, 8'sb11111111, 8'sb00001101, 8'sb00000000, 8'sb11110011, 8'sb11111101, 8'sb11110111, 8'sb11100100, 8'sb00001010, 8'sb00011111, 8'sb11101110, 8'sb11011011, 8'sb11100101, 8'sb11110100, 8'sb11111101, 8'sb00001110, 8'sb00000110, 8'sb11110111, 8'sb11101010, 8'sb11101001, 8'sb11110011, 8'sb11101000, 8'sb00010011, 8'sb00010100, 8'sb11011000, 8'sb00010110, 8'sb11110001, 8'sb11110110, 8'sb11101110, 8'sb00010101, 8'sb00001101, 8'sb11100010, 8'sb11110001, 8'sb11101110, 8'sb11110111, 8'sb11111100, 8'sb00000100, 8'sb11111011, 8'sb11110010, 8'sb11110010, 8'sb00010000, 8'sb00001101, 8'sb11111011, 8'sb11111001, 8'sb11100001, 8'sb11010011, 8'sb00001000, 8'sb00000110, 8'sb00000111, 8'sb00001000, 8'sb00000100, 8'sb11101101, 8'sb00001011, 8'sb00000100, 8'sb00100000, 8'sb00001101, 8'sb11111001, 8'sb11111001, 8'sb11110110, 8'sb00001111, 8'sb00000110, 8'sb00010111, 8'sb00100000, 8'sb00011110, 8'sb11111001, 8'sb11111101, 8'sb11101110, 8'sb00010010, 8'sb11110011, 8'sb00010110, 8'sb00010111, 8'sb00101010, 8'sb00110110, 8'sb00101010, 8'sb00110000, 8'sb00001111, 8'sb00011111, 8'sb00111101, 8'sb00001110, 8'sb11100100, 8'sb11110101, 8'sb11111010, 8'sb11101010, 8'sb00000000, 8'sb00011111, 8'sb00011011, 8'sb00100011, 8'sb00111000, 8'sb00101001, 8'sb00101101, 8'sb00010100, 8'sb00011110, 8'sb00101010, 8'sb00000011, 8'sb00001001, 8'sb00000100, 8'sb00000100, 8'sb11110001, 8'sb11100000, 8'sb00010001, 8'sb00010010, 8'sb11110000, 8'sb11101101, 8'sb11111110, 8'sb00001001, 8'sb00000101, 8'sb00001010, 8'sb11111110,
    8'sb00001100, 8'sb00000010, 8'sb11111000, 8'sb11011100, 8'sb11100010, 8'sb11101000, 8'sb11110010, 8'sb11111010, 8'sb10111001, 8'sb11001100, 8'sb11010110, 8'sb11101001, 8'sb11110100, 8'sb00000101, 8'sb00000010, 8'sb11010110, 8'sb11010001, 8'sb11010111, 8'sb10110011, 8'sb11000000, 8'sb10111011, 8'sb11010100, 8'sb11011101, 8'sb10111111, 8'sb11100010, 8'sb11111011, 8'sb11110000, 8'sb11100101, 8'sb11110101, 8'sb00001000, 8'sb00000010, 8'sb00001010, 8'sb11101101, 8'sb11101101, 8'sb00000101, 8'sb00000100, 8'sb00000000, 8'sb00001101, 8'sb00010110, 8'sb00001111, 8'sb11110100, 8'sb11011111, 8'sb00001101, 8'sb00101000, 8'sb00110010, 8'sb00001100, 8'sb11110110, 8'sb11110010, 8'sb11101001, 8'sb11101000, 8'sb11011111, 8'sb11111111, 8'sb11111100, 8'sb00110100, 8'sb00011000, 8'sb00000001, 8'sb00100011, 8'sb00101010, 8'sb00010001, 8'sb00000101, 8'sb00001010, 8'sb11110010, 8'sb00000011, 8'sb11111001, 8'sb00000001, 8'sb00100001, 8'sb00101000, 8'sb00101110, 8'sb00010010, 8'sb00000100, 8'sb00110110, 8'sb00010010, 8'sb11101100, 8'sb11110011, 8'sb00000101, 8'sb00010011, 8'sb00011000, 8'sb11111101, 8'sb00000001, 8'sb00001111, 8'sb00001011, 8'sb00011001, 8'sb11100011, 8'sb11100010, 8'sb00100101, 8'sb11110111, 8'sb11100100, 8'sb00001100, 8'sb00100001, 8'sb00100000, 8'sb00000001, 8'sb11101010, 8'sb11111110, 8'sb11110110, 8'sb00000001, 8'sb00001001, 8'sb00011010, 8'sb11100101, 8'sb11111100, 8'sb00000011, 8'sb00000110, 8'sb00010110, 8'sb00100010, 8'sb00001010, 8'sb11101000, 8'sb00000000, 8'sb00011000, 8'sb00011100, 8'sb11111001, 8'sb00001011, 8'sb00000001, 8'sb00000101, 8'sb00000000, 8'sb11101100, 8'sb11111010, 8'sb00110101, 8'sb00110000, 8'sb11101100, 8'sb11110101, 8'sb00100101, 8'sb00011011, 8'sb00000111, 8'sb00010111, 8'sb00010001, 8'sb11111001, 8'sb11111000, 8'sb11100011, 8'sb00000011, 8'sb00000111, 8'sb00011000, 8'sb00011011, 8'sb11010000, 8'sb11100110, 8'sb00001101, 8'sb00000010, 8'sb11110010, 8'sb11111011, 8'sb00000001, 8'sb11111011, 8'sb00000010, 8'sb00010011, 8'sb00010000, 8'sb00000011, 8'sb00001111, 8'sb00000001, 8'sb11011011, 8'sb11110001, 8'sb11111101, 8'sb11111011, 8'sb11111111, 8'sb11111011, 8'sb11101101, 8'sb11001010, 8'sb00001001, 8'sb11111000, 8'sb11010010, 8'sb11111101, 8'sb00100011, 8'sb00001001, 8'sb00001000, 8'sb11111101, 8'sb00000011, 8'sb00001011, 8'sb00010110, 8'sb00001000, 8'sb11111110, 8'sb11010001, 8'sb11101111, 8'sb00001011, 8'sb11011110, 8'sb11100111, 8'sb11100111, 8'sb11101110, 8'sb00000010, 8'sb11111111, 8'sb11111000, 8'sb11110100, 8'sb11101100, 8'sb11101010, 8'sb11011111, 8'sb11001010, 8'sb00000011, 8'sb00001000, 8'sb11110001, 8'sb11100101, 8'sb11010110, 8'sb11010011, 8'sb11001100, 8'sb11001001, 8'sb10110111, 8'sb11000101, 8'sb10110101, 8'sb10101001, 8'sb11100000, 8'sb11100111, 8'sb11111111,
    8'sb11110100, 8'sb00000000, 8'sb00000000, 8'sb11111011, 8'sb11111010, 8'sb11101000, 8'sb11110001, 8'sb00001011, 8'sb11101110, 8'sb00011010, 8'sb00011110, 8'sb00000001, 8'sb00001100, 8'sb00000011, 8'sb00000101, 8'sb11110010, 8'sb11110110, 8'sb11111001, 8'sb00010000, 8'sb11101111, 8'sb00000011, 8'sb00000011, 8'sb11110011, 8'sb11101101, 8'sb00000100, 8'sb00000001, 8'sb11111111, 8'sb11101111, 8'sb00001000, 8'sb00001100, 8'sb11101011, 8'sb11011000, 8'sb11010010, 8'sb11011100, 8'sb11101110, 8'sb11101111, 8'sb11111101, 8'sb00001010, 8'sb00001110, 8'sb00010101, 8'sb00001101, 8'sb11111001, 8'sb11100110, 8'sb11101001, 8'sb10111100, 8'sb10111001, 8'sb10111011, 8'sb11010111, 8'sb11110101, 8'sb00001100, 8'sb00000000, 8'sb00010010, 8'sb00100101, 8'sb00001011, 8'sb00010110, 8'sb00100000, 8'sb11011010, 8'sb11001011, 8'sb11001100, 8'sb11001011, 8'sb11001010, 8'sb11111100, 8'sb00011001, 8'sb00001100, 8'sb11101100, 8'sb11111001, 8'sb11111011, 8'sb11110101, 8'sb00010110, 8'sb11111101, 8'sb11010101, 8'sb11011001, 8'sb11100110, 8'sb11011010, 8'sb11110101, 8'sb00100001, 8'sb00001100, 8'sb11111111, 8'sb11100010, 8'sb11010100, 8'sb11100010, 8'sb11010010, 8'sb11100000, 8'sb11011111, 8'sb11101111, 8'sb11110101, 8'sb00001000, 8'sb00001001, 8'sb00000101, 8'sb00000010, 8'sb11111001, 8'sb00011000, 8'sb00000000, 8'sb11110011, 8'sb00000101, 8'sb11010000, 8'sb11001110, 8'sb11101101, 8'sb11101111, 8'sb00101000, 8'sb00010001, 8'sb00011011, 8'sb00010001, 8'sb11111010, 8'sb00010001, 8'sb00011001, 8'sb00011000, 8'sb11100001, 8'sb11010101, 8'sb11011001, 8'sb11111000, 8'sb01000001, 8'sb11101010, 8'sb00100000, 8'sb00000111, 8'sb00100001, 8'sb00011101, 8'sb00010110, 8'sb00010001, 8'sb00101001, 8'sb11101011, 8'sb11011001, 8'sb11110000, 8'sb11101000, 8'sb11111011, 8'sb01011110, 8'sb11101100, 8'sb00000100, 8'sb11101100, 8'sb11111101, 8'sb00011000, 8'sb00000100, 8'sb00001111, 8'sb00010010, 8'sb11110100, 8'sb11111011, 8'sb00001001, 8'sb00010000, 8'sb01000001, 8'sb00111101, 8'sb11111011, 8'sb11101111, 8'sb00001010, 8'sb11110110, 8'sb11111011, 8'sb11110101, 8'sb11101001, 8'sb00001011, 8'sb00101101, 8'sb00101101, 8'sb00110101, 8'sb00011101, 8'sb00111110, 8'sb00000001, 8'sb00010110, 8'sb11110110, 8'sb00100000, 8'sb11111100, 8'sb11111001, 8'sb11111011, 8'sb11110101, 8'sb11110011, 8'sb00001111, 8'sb00110011, 8'sb00110101, 8'sb00100100, 8'sb11111011, 8'sb11111110, 8'sb00000011, 8'sb11010000, 8'sb11000101, 8'sb11100100, 8'sb11101111, 8'sb11101011, 8'sb11100110, 8'sb11100000, 8'sb11001110, 8'sb11100110, 8'sb00010011, 8'sb00011011, 8'sb00001000, 8'sb00010111, 8'sb00000111, 8'sb00001010, 8'sb00001010, 8'sb00011011, 8'sb00001001, 8'sb00001101, 8'sb00100001, 8'sb00000111, 8'sb11111110, 8'sb11001011, 8'sb11111000, 8'sb11110011, 8'sb00000101, 8'sb00001100,
    8'sb00001001, 8'sb00000110, 8'sb11111110, 8'sb00011101, 8'sb00011111, 8'sb11111000, 8'sb00000001, 8'sb11011010, 8'sb00000010, 8'sb00111110, 8'sb00111111, 8'sb00100101, 8'sb11111001, 8'sb11110111, 8'sb11110101, 8'sb11110011, 8'sb00010100, 8'sb00101100, 8'sb00101100, 8'sb00101010, 8'sb00001011, 8'sb11111110, 8'sb00010100, 8'sb00001011, 8'sb00000100, 8'sb00010001, 8'sb11111110, 8'sb11111000, 8'sb00000110, 8'sb11101000, 8'sb00000111, 8'sb11111111, 8'sb00010101, 8'sb00000010, 8'sb11111010, 8'sb11011011, 8'sb11110110, 8'sb11111100, 8'sb11110011, 8'sb11100000, 8'sb11101111, 8'sb11110100, 8'sb11100011, 8'sb00001110, 8'sb00010100, 8'sb00010110, 8'sb00011000, 8'sb00000010, 8'sb00000010, 8'sb00001011, 8'sb00000001, 8'sb11011111, 8'sb11100101, 8'sb11100000, 8'sb00001001, 8'sb11111000, 8'sb11110101, 8'sb00000011, 8'sb00100110, 8'sb00000011, 8'sb11110110, 8'sb11110010, 8'sb11101011, 8'sb11111110, 8'sb11110001, 8'sb11011011, 8'sb11111001, 8'sb11111001, 8'sb11101001, 8'sb11111110, 8'sb11011100, 8'sb00000111, 8'sb00001011, 8'sb00001010, 8'sb00000010, 8'sb11101101, 8'sb11010100, 8'sb11010011, 8'sb11111001, 8'sb00000100, 8'sb00001001, 8'sb00000001, 8'sb11011100, 8'sb11000110, 8'sb11111100, 8'sb11110000, 8'sb00001011, 8'sb00001011, 8'sb00000011, 8'sb11110011, 8'sb11101001, 8'sb11111110, 8'sb00000111, 8'sb00001010, 8'sb00011001, 8'sb00010101, 8'sb00010111, 8'sb11111010, 8'sb11100001, 8'sb00010111, 8'sb11111011, 8'sb00010010, 8'sb00000110, 8'sb00011011, 8'sb00100011, 8'sb00010110, 8'sb00100011, 8'sb00101011, 8'sb00101100, 8'sb00010011, 8'sb11110100, 8'sb01001010, 8'sb11110100, 8'sb00000110, 8'sb11111011, 8'sb00011100, 8'sb00001101, 8'sb00011100, 8'sb00011101, 8'sb00010111, 8'sb00101100, 8'sb00100000, 8'sb00011011, 8'sb00000101, 8'sb11111010, 8'sb00101010, 8'sb11010110, 8'sb00000101, 8'sb00010010, 8'sb00001110, 8'sb11110001, 8'sb11110111, 8'sb11111100, 8'sb00010010, 8'sb00100011, 8'sb00001010, 8'sb00000011, 8'sb11110000, 8'sb11111011, 8'sb00110111, 8'sb11110111, 8'sb00011011, 8'sb11111000, 8'sb11111001, 8'sb11101011, 8'sb11101111, 8'sb11111011, 8'sb00010000, 8'sb11111111, 8'sb11110110, 8'sb11010001, 8'sb11011000, 8'sb11111101, 8'sb11110000, 8'sb11111110, 8'sb00000100, 8'sb11100011, 8'sb11101001, 8'sb11110101, 8'sb00000111, 8'sb11110000, 8'sb11101011, 8'sb11010001, 8'sb11000101, 8'sb11110001, 8'sb11101010, 8'sb11111110, 8'sb11100011, 8'sb00000111, 8'sb11100010, 8'sb11110000, 8'sb00010000, 8'sb00011000, 8'sb00010001, 8'sb11110001, 8'sb00010110, 8'sb11101101, 8'sb11011100, 8'sb00010000, 8'sb11110100, 8'sb11110110, 8'sb00001101, 8'sb00001000, 8'sb00001110, 8'sb00110100, 8'sb00111001, 8'sb00101101, 8'sb00011110, 8'sb00011001, 8'sb00100111, 8'sb11111001, 8'sb11101011, 8'sb00000110, 8'sb11110100, 8'sb00001010, 8'sb11111011,
    8'sb00001010, 8'sb00000110, 8'sb00001010, 8'sb00000111, 8'sb00010100, 8'sb00010111, 8'sb00100011, 8'sb00010111, 8'sb00100110, 8'sb00101111, 8'sb00100010, 8'sb00000111, 8'sb11110111, 8'sb00000110, 8'sb00000000, 8'sb00010100, 8'sb11111001, 8'sb00001100, 8'sb11110111, 8'sb11101001, 8'sb11011101, 8'sb11100111, 8'sb00010111, 8'sb00111011, 8'sb00101110, 8'sb01000001, 8'sb00010001, 8'sb00010100, 8'sb00000110, 8'sb11101111, 8'sb11011010, 8'sb11010011, 8'sb11011111, 8'sb11010100, 8'sb11010000, 8'sb11100111, 8'sb00010010, 8'sb00101001, 8'sb00010011, 8'sb00000001, 8'sb00011010, 8'sb00101111, 8'sb11101011, 8'sb11110010, 8'sb11100000, 8'sb11011100, 8'sb11101010, 8'sb11111101, 8'sb11111000, 8'sb00000111, 8'sb00011110, 8'sb00110101, 8'sb00101110, 8'sb00100101, 8'sb00010011, 8'sb00000110, 8'sb11101110, 8'sb11111000, 8'sb11011111, 8'sb11100111, 8'sb11101110, 8'sb00000111, 8'sb00101000, 8'sb00010100, 8'sb00001010, 8'sb00000110, 8'sb00001110, 8'sb00000110, 8'sb00011101, 8'sb11111010, 8'sb11111010, 8'sb11110001, 8'sb11100001, 8'sb00000010, 8'sb11111010, 8'sb00001010, 8'sb00010110, 8'sb11110101, 8'sb11010011, 8'sb11011101, 8'sb11100010, 8'sb11111011, 8'sb00100001, 8'sb00000001, 8'sb00100001, 8'sb00000110, 8'sb11010111, 8'sb11111101, 8'sb11111001, 8'sb00000010, 8'sb00010011, 8'sb11101110, 8'sb11101001, 8'sb11100110, 8'sb11011010, 8'sb00000001, 8'sb00001001, 8'sb00000101, 8'sb00010111, 8'sb11010001, 8'sb11110001, 8'sb11111100, 8'sb00001001, 8'sb00000110, 8'sb00001101, 8'sb11110101, 8'sb11101110, 8'sb11101010, 8'sb11110000, 8'sb11011111, 8'sb00000101, 8'sb11010010, 8'sb11110000, 8'sb11101100, 8'sb11101010, 8'sb11111011, 8'sb00011101, 8'sb00000110, 8'sb11101101, 8'sb11110000, 8'sb00000100, 8'sb11101111, 8'sb11111111, 8'sb11101001, 8'sb11011111, 8'sb11011010, 8'sb00011110, 8'sb11001010, 8'sb00000010, 8'sb00001101, 8'sb00011010, 8'sb11111010, 8'sb11001101, 8'sb11110011, 8'sb00000011, 8'sb11111011, 8'sb11111010, 8'sb11101101, 8'sb11100001, 8'sb11101100, 8'sb00000011, 8'sb11011000, 8'sb00000000, 8'sb00011010, 8'sb00010111, 8'sb00011001, 8'sb00001001, 8'sb11110010, 8'sb11111011, 8'sb00000100, 8'sb11111111, 8'sb11110011, 8'sb11100100, 8'sb11101001, 8'sb11110111, 8'sb00000010, 8'sb11111111, 8'sb00001100, 8'sb00010100, 8'sb00011101, 8'sb00100101, 8'sb00010001, 8'sb00000011, 8'sb11110110, 8'sb11101010, 8'sb11111110, 8'sb00000110, 8'sb11100101, 8'sb11111101, 8'sb11110110, 8'sb11101010, 8'sb00000011, 8'sb00010111, 8'sb00100110, 8'sb00101110, 8'sb00110000, 8'sb00100110, 8'sb00100111, 8'sb00001000, 8'sb11111110, 8'sb11110011, 8'sb11101110, 8'sb00000101, 8'sb00000100, 8'sb11100100, 8'sb11011101, 8'sb11101010, 8'sb00000110, 8'sb00101100, 8'sb11110100, 8'sb00010101, 8'sb00000011, 8'sb11111100, 8'sb00011111, 8'sb00001001, 8'sb00001100,
    8'sb00001000, 8'sb11111100, 8'sb11110110, 8'sb11100001, 8'sb11100100, 8'sb11011101, 8'sb11100010, 8'sb11100111, 8'sb11011010, 8'sb11100110, 8'sb11101010, 8'sb11100010, 8'sb11110111, 8'sb00000100, 8'sb00000000, 8'sb11101001, 8'sb11010101, 8'sb11011001, 8'sb10110011, 8'sb10011011, 8'sb10011101, 8'sb10111001, 8'sb11011101, 8'sb00000011, 8'sb11111111, 8'sb11110011, 8'sb00001000, 8'sb00000100, 8'sb11110101, 8'sb11001000, 8'sb11010110, 8'sb11101000, 8'sb11100101, 8'sb11101001, 8'sb11110010, 8'sb11110100, 8'sb11111010, 8'sb11111011, 8'sb11111111, 8'sb00001001, 8'sb00100000, 8'sb00001010, 8'sb11111010, 8'sb00000101, 8'sb11111101, 8'sb00001011, 8'sb00001011, 8'sb00001000, 8'sb00000000, 8'sb00000010, 8'sb00010111, 8'sb00011010, 8'sb00010110, 8'sb00010101, 8'sb00011111, 8'sb00011110, 8'sb00010010, 8'sb11111111, 8'sb00010111, 8'sb00100011, 8'sb00101010, 8'sb00010000, 8'sb11111010, 8'sb11111011, 8'sb00000111, 8'sb00011000, 8'sb00001001, 8'sb00010000, 8'sb01010010, 8'sb01010010, 8'sb00010101, 8'sb00000100, 8'sb00100110, 8'sb00111011, 8'sb00101000, 8'sb00100111, 8'sb00011100, 8'sb11100110, 8'sb11100000, 8'sb00000010, 8'sb00000101, 8'sb00010110, 8'sb00111000, 8'sb01011101, 8'sb00110011, 8'sb00011010, 8'sb00110110, 8'sb00101000, 8'sb00011111, 8'sb00101001, 8'sb00000100, 8'sb11111110, 8'sb11110010, 8'sb11111111, 8'sb00011110, 8'sb11111010, 8'sb11111101, 8'sb00110101, 8'sb00011111, 8'sb00000001, 8'sb11101110, 8'sb11101111, 8'sb00001011, 8'sb00010101, 8'sb00001110, 8'sb00000010, 8'sb11111110, 8'sb11111110, 8'sb11111000, 8'sb00000001, 8'sb11101110, 8'sb11001010, 8'sb11011101, 8'sb11111100, 8'sb11010011, 8'sb11011110, 8'sb11101001, 8'sb11110101, 8'sb00011000, 8'sb00001101, 8'sb00000110, 8'sb11110000, 8'sb11110011, 8'sb00000101, 8'sb11111100, 8'sb11011100, 8'sb00011010, 8'sb11011011, 8'sb11110101, 8'sb11101101, 8'sb11011101, 8'sb11100101, 8'sb11110100, 8'sb00000100, 8'sb11110101, 8'sb11100010, 8'sb11110010, 8'sb00000000, 8'sb00000100, 8'sb11101100, 8'sb11101011, 8'sb10101100, 8'sb11110110, 8'sb11111101, 8'sb11110100, 8'sb11100001, 8'sb00000111, 8'sb11110100, 8'sb11110100, 8'sb11110000, 8'sb11111000, 8'sb00010101, 8'sb00001110, 8'sb11001010, 8'sb11110001, 8'sb11010110, 8'sb11110010, 8'sb00010011, 8'sb00001001, 8'sb00001010, 8'sb11111010, 8'sb00000010, 8'sb11111010, 8'sb11101000, 8'sb00000001, 8'sb00001000, 8'sb00011110, 8'sb00001110, 8'sb11110100, 8'sb00010010, 8'sb11111100, 8'sb11101101, 8'sb00001011, 8'sb00011100, 8'sb00011110, 8'sb00100110, 8'sb00010000, 8'sb00001001, 8'sb00000100, 8'sb00010010, 8'sb11101100, 8'sb11100110, 8'sb11110100, 8'sb11111101, 8'sb11001001, 8'sb11100010, 8'sb00000111, 8'sb00001111, 8'sb00100000, 8'sb00010000, 8'sb00011011, 8'sb00010010, 8'sb11111110, 8'sb00010100, 8'sb11101100, 8'sb11111010,
    8'sb00000110, 8'sb11111110, 8'sb00000111, 8'sb00001100, 8'sb00001000, 8'sb00100010, 8'sb00011011, 8'sb00100111, 8'sb00100111, 8'sb00011111, 8'sb00100010, 8'sb00010001, 8'sb11111100, 8'sb11111100, 8'sb00001100, 8'sb00001111, 8'sb00000100, 8'sb11111101, 8'sb11111010, 8'sb11011110, 8'sb11111111, 8'sb11111110, 8'sb00011011, 8'sb11110000, 8'sb11101110, 8'sb11101110, 8'sb00001011, 8'sb11100010, 8'sb00000011, 8'sb00000111, 8'sb11001111, 8'sb11100001, 8'sb11100001, 8'sb11100101, 8'sb11111100, 8'sb00000111, 8'sb00001000, 8'sb00001100, 8'sb00100001, 8'sb11110110, 8'sb11101000, 8'sb00011000, 8'sb11011111, 8'sb11100011, 8'sb10100010, 8'sb11001000, 8'sb11011101, 8'sb11111000, 8'sb00000100, 8'sb00001110, 8'sb00010101, 8'sb00011010, 8'sb00010000, 8'sb00000110, 8'sb11110011, 8'sb11011000, 8'sb11011111, 8'sb11011101, 8'sb11000111, 8'sb11111110, 8'sb00000010, 8'sb00000100, 8'sb00001000, 8'sb00100010, 8'sb00011000, 8'sb00001000, 8'sb00001110, 8'sb00000011, 8'sb00000000, 8'sb11111010, 8'sb11101111, 8'sb11011111, 8'sb11111001, 8'sb00010001, 8'sb00001001, 8'sb11111010, 8'sb00000011, 8'sb00011011, 8'sb00001010, 8'sb00001100, 8'sb00010111, 8'sb00100100, 8'sb00011000, 8'sb00001011, 8'sb11011001, 8'sb11110111, 8'sb00011010, 8'sb00010000, 8'sb11111111, 8'sb11010010, 8'sb00000010, 8'sb00100000, 8'sb11110111, 8'sb00001001, 8'sb00010010, 8'sb00110110, 8'sb00010001, 8'sb11111001, 8'sb11011111, 8'sb11110110, 8'sb00000111, 8'sb11111010, 8'sb11111001, 8'sb11111000, 8'sb00101010, 8'sb00001010, 8'sb11101110, 8'sb11110010, 8'sb11101111, 8'sb11101010, 8'sb11110111, 8'sb11110111, 8'sb00011111, 8'sb11110011, 8'sb00001100, 8'sb00001001, 8'sb00010000, 8'sb00011000, 8'sb00001011, 8'sb11101111, 8'sb11100010, 8'sb11100100, 8'sb11010100, 8'sb11100011, 8'sb11110000, 8'sb11101001, 8'sb00000110, 8'sb11011000, 8'sb11110100, 8'sb00001010, 8'sb00010110, 8'sb00010011, 8'sb11111010, 8'sb11110111, 8'sb11110001, 8'sb11111001, 8'sb11110101, 8'sb00010110, 8'sb00011011, 8'sb11101110, 8'sb00010111, 8'sb11111110, 8'sb00100010, 8'sb00101101, 8'sb00011110, 8'sb00000000, 8'sb00000011, 8'sb00001110, 8'sb00010001, 8'sb00010001, 8'sb00000010, 8'sb00010011, 8'sb00101010, 8'sb00000011, 8'sb00010110, 8'sb11111001, 8'sb00000101, 8'sb00010111, 8'sb00011000, 8'sb00001000, 8'sb00001110, 8'sb00000111, 8'sb00000011, 8'sb11101001, 8'sb11110001, 8'sb00001110, 8'sb00011010, 8'sb11110011, 8'sb11111111, 8'sb11101110, 8'sb11011000, 8'sb11100111, 8'sb00000010, 8'sb00000010, 8'sb00000000, 8'sb11111100, 8'sb00001101, 8'sb00001010, 8'sb00001110, 8'sb00001010, 8'sb00010000, 8'sb11111001, 8'sb11111010, 8'sb00011001, 8'sb00011110, 8'sb00011011, 8'sb00010010, 8'sb00010110, 8'sb00010010, 8'sb00011111, 8'sb00010100, 8'sb00011010, 8'sb00011110, 8'sb11111111, 8'sb00011000, 8'sb00000111,
    8'sb11111111, 8'sb11110110, 8'sb00001000, 8'sb00011011, 8'sb00001000, 8'sb00011001, 8'sb00001001, 8'sb11111000, 8'sb00011000, 8'sb00011101, 8'sb00101111, 8'sb00011111, 8'sb11110100, 8'sb00000011, 8'sb11111101, 8'sb00011100, 8'sb00010100, 8'sb11111111, 8'sb00011011, 8'sb00001001, 8'sb11101110, 8'sb11101010, 8'sb00001010, 8'sb00011011, 8'sb00000010, 8'sb00001000, 8'sb00001110, 8'sb00010001, 8'sb11110111, 8'sb00001011, 8'sb11101111, 8'sb11101100, 8'sb11110100, 8'sb00010010, 8'sb00010001, 8'sb11110111, 8'sb00001100, 8'sb00010001, 8'sb00000011, 8'sb11111110, 8'sb00001000, 8'sb00001101, 8'sb11011111, 8'sb11100001, 8'sb11100011, 8'sb11110111, 8'sb00010100, 8'sb00010111, 8'sb00010001, 8'sb00001001, 8'sb00001100, 8'sb00010011, 8'sb00001010, 8'sb00001001, 8'sb00011101, 8'sb00100111, 8'sb11110000, 8'sb11001101, 8'sb11110101, 8'sb00000100, 8'sb11111101, 8'sb00001010, 8'sb11110010, 8'sb11011000, 8'sb11001100, 8'sb11100010, 8'sb11101011, 8'sb11110010, 8'sb11100010, 8'sb00000110, 8'sb11010010, 8'sb11001111, 8'sb00000100, 8'sb00001000, 8'sb11111101, 8'sb00001000, 8'sb11100110, 8'sb11011011, 8'sb11111001, 8'sb11101101, 8'sb11010000, 8'sb10101111, 8'sb11001110, 8'sb00001110, 8'sb11100111, 8'sb11100011, 8'sb11101000, 8'sb11110000, 8'sb00000111, 8'sb00010010, 8'sb00001011, 8'sb00000110, 8'sb00000110, 8'sb00010111, 8'sb00001101, 8'sb11100100, 8'sb11011110, 8'sb00101010, 8'sb11100111, 8'sb00010110, 8'sb11111100, 8'sb00001011, 8'sb11111111, 8'sb00000001, 8'sb11110110, 8'sb00000101, 8'sb00010111, 8'sb00000111, 8'sb11110111, 8'sb11110001, 8'sb00001011, 8'sb00110001, 8'sb11011111, 8'sb00100011, 8'sb11111001, 8'sb11111111, 8'sb11110000, 8'sb11101000, 8'sb11111100, 8'sb00011000, 8'sb00100011, 8'sb00011100, 8'sb00001110, 8'sb00000111, 8'sb00101010, 8'sb00011111, 8'sb11100100, 8'sb00100000, 8'sb00010011, 8'sb00000001, 8'sb00000011, 8'sb11111011, 8'sb11110110, 8'sb00010010, 8'sb00010101, 8'sb00001101, 8'sb00001000, 8'sb00001001, 8'sb00101001, 8'sb00100011, 8'sb11111010, 8'sb00100110, 8'sb00100001, 8'sb00010001, 8'sb00010111, 8'sb11111110, 8'sb11111111, 8'sb00000101, 8'sb00000000, 8'sb00001101, 8'sb00010010, 8'sb00011011, 8'sb00100100, 8'sb11101101, 8'sb11111111, 8'sb00011111, 8'sb00010110, 8'sb00000010, 8'sb00001011, 8'sb00000111, 8'sb11110011, 8'sb11110001, 8'sb11111000, 8'sb00001011, 8'sb00001110, 8'sb00010111, 8'sb00110010, 8'sb00001101, 8'sb00001011, 8'sb11101011, 8'sb11100101, 8'sb00001011, 8'sb00000101, 8'sb11110011, 8'sb11110000, 8'sb11110010, 8'sb00000100, 8'sb00010111, 8'sb00101110, 8'sb01000100, 8'sb00110111, 8'sb11111000, 8'sb00001000, 8'sb00000000, 8'sb11101101, 8'sb11110001, 8'sb11110001, 8'sb00001111, 8'sb11111010, 8'sb00010001, 8'sb11110101, 8'sb11011010, 8'sb00010111, 8'sb00010000, 8'sb11111111, 8'sb11111000,
    8'sb11111111, 8'sb00000010, 8'sb11111100, 8'sb11101001, 8'sb11100100, 8'sb11011100, 8'sb11010011, 8'sb11011001, 8'sb11010101, 8'sb11010011, 8'sb11010111, 8'sb11101001, 8'sb11110100, 8'sb11110110, 8'sb11111011, 8'sb11100010, 8'sb00001001, 8'sb11011101, 8'sb10111011, 8'sb11011101, 8'sb11001101, 8'sb11011001, 8'sb11111010, 8'sb00001100, 8'sb00010111, 8'sb11110010, 8'sb00000001, 8'sb11111000, 8'sb00000000, 8'sb00001101, 8'sb11110001, 8'sb11100001, 8'sb11000011, 8'sb11100110, 8'sb11111001, 8'sb00000000, 8'sb00001010, 8'sb00001011, 8'sb00011101, 8'sb00010110, 8'sb00100010, 8'sb11110101, 8'sb11100011, 8'sb11110001, 8'sb11101011, 8'sb11011011, 8'sb11100101, 8'sb11111110, 8'sb00010100, 8'sb00011000, 8'sb00010110, 8'sb00100000, 8'sb00011110, 8'sb00010011, 8'sb00011000, 8'sb00011001, 8'sb11001011, 8'sb11110100, 8'sb11101010, 8'sb11100110, 8'sb11111110, 8'sb00000010, 8'sb00001000, 8'sb00001101, 8'sb00010110, 8'sb00010110, 8'sb00001000, 8'sb00001110, 8'sb00100110, 8'sb00011101, 8'sb11000010, 8'sb11011011, 8'sb11110001, 8'sb11110001, 8'sb00000111, 8'sb11111000, 8'sb11110110, 8'sb11111011, 8'sb00010110, 8'sb00001000, 8'sb11100110, 8'sb11110011, 8'sb00100101, 8'sb00010000, 8'sb11100000, 8'sb11110010, 8'sb11111011, 8'sb00000101, 8'sb11111011, 8'sb00000100, 8'sb00010110, 8'sb00100110, 8'sb00100000, 8'sb00010011, 8'sb11110000, 8'sb11100001, 8'sb11001010, 8'sb11110000, 8'sb11110101, 8'sb11111110, 8'sb00001100, 8'sb11111110, 8'sb00000011, 8'sb11111011, 8'sb00010011, 8'sb00010000, 8'sb00010111, 8'sb11111000, 8'sb11101001, 8'sb11100000, 8'sb11010111, 8'sb11011010, 8'sb00001110, 8'sb11110001, 8'sb11110110, 8'sb11111110, 8'sb11111110, 8'sb11111111, 8'sb00001110, 8'sb00010011, 8'sb00010111, 8'sb00000110, 8'sb11101111, 8'sb11001111, 8'sb11001010, 8'sb11010101, 8'sb11101011, 8'sb00010011, 8'sb00011001, 8'sb11111111, 8'sb11111001, 8'sb11111101, 8'sb00000010, 8'sb00100000, 8'sb00010000, 8'sb00000101, 8'sb11110000, 8'sb10101000, 8'sb10100111, 8'sb11111110, 8'sb11110111, 8'sb00000001, 8'sb00001100, 8'sb11111111, 8'sb11111001, 8'sb11101110, 8'sb11101100, 8'sb00000010, 8'sb00000110, 8'sb11111111, 8'sb11011001, 8'sb10111011, 8'sb10111100, 8'sb11101010, 8'sb00001000, 8'sb00001101, 8'sb00000001, 8'sb11110110, 8'sb00000011, 8'sb00011011, 8'sb00001001, 8'sb11111011, 8'sb11111001, 8'sb11111011, 8'sb00010001, 8'sb11110010, 8'sb11101000, 8'sb11111100, 8'sb11110110, 8'sb00111111, 8'sb00101100, 8'sb00101110, 8'sb00100101, 8'sb00011101, 8'sb00010001, 8'sb00000100, 8'sb00000001, 8'sb00001110, 8'sb00110000, 8'sb00101011, 8'sb11100101, 8'sb11101111, 8'sb00001010, 8'sb00001100, 8'sb00101101, 8'sb00010111, 8'sb11111111, 8'sb00010110, 8'sb00010100, 8'sb00000100, 8'sb11110110, 8'sb11100001, 8'sb00010011, 8'sb00000000, 8'sb00100011, 8'sb00000111,
    8'sb00000101, 8'sb11111111, 8'sb00000100, 8'sb00011011, 8'sb00101001, 8'sb00110110, 8'sb01000111, 8'sb00011010, 8'sb00010111, 8'sb00111101, 8'sb00101011, 8'sb00100100, 8'sb11111001, 8'sb00001010, 8'sb00001001, 8'sb00100101, 8'sb00110111, 8'sb00100110, 8'sb00101110, 8'sb00110010, 8'sb00111000, 8'sb01000110, 8'sb00100110, 8'sb00110111, 8'sb00101100, 8'sb00001110, 8'sb11101011, 8'sb11101001, 8'sb11111110, 8'sb00100010, 8'sb00111001, 8'sb00011010, 8'sb00011110, 8'sb00001101, 8'sb00001100, 8'sb00010010, 8'sb00011101, 8'sb00011001, 8'sb00011011, 8'sb00011000, 8'sb00001001, 8'sb00101100, 8'sb00001111, 8'sb11111010, 8'sb00011100, 8'sb00000110, 8'sb00000110, 8'sb11101110, 8'sb11101011, 8'sb11110110, 8'sb11100001, 8'sb11110010, 8'sb11110111, 8'sb00001001, 8'sb00100011, 8'sb00011000, 8'sb11011100, 8'sb11110001, 8'sb00001111, 8'sb00001000, 8'sb11111100, 8'sb11111010, 8'sb00000010, 8'sb11110010, 8'sb11011110, 8'sb11100101, 8'sb11101101, 8'sb11110111, 8'sb11011111, 8'sb00010100, 8'sb11011100, 8'sb00000110, 8'sb00001001, 8'sb11111100, 8'sb11101100, 8'sb11111111, 8'sb00100110, 8'sb00010111, 8'sb11110111, 8'sb11111011, 8'sb11110100, 8'sb11101001, 8'sb11111010, 8'sb00011000, 8'sb11001001, 8'sb11100010, 8'sb11101001, 8'sb11011110, 8'sb00000001, 8'sb11111110, 8'sb00100010, 8'sb00011101, 8'sb00011001, 8'sb00000110, 8'sb11100011, 8'sb11111011, 8'sb11010101, 8'sb11110110, 8'sb00000100, 8'sb00000111, 8'sb11010000, 8'sb11110111, 8'sb11110100, 8'sb11011111, 8'sb00001110, 8'sb00110000, 8'sb00000111, 8'sb11110011, 8'sb11101101, 8'sb11111010, 8'sb00001100, 8'sb11101001, 8'sb00100110, 8'sb00111001, 8'sb11111011, 8'sb11101100, 8'sb11011110, 8'sb11010100, 8'sb00010011, 8'sb00001010, 8'sb11100101, 8'sb00000100, 8'sb00001111, 8'sb00011010, 8'sb00010000, 8'sb11101000, 8'sb11011101, 8'sb00101101, 8'sb00011100, 8'sb00000101, 8'sb11111001, 8'sb11100001, 8'sb11111011, 8'sb00001000, 8'sb00100000, 8'sb00001101, 8'sb00010010, 8'sb00001010, 8'sb11110010, 8'sb11110101, 8'sb00010010, 8'sb00011110, 8'sb11111100, 8'sb00011101, 8'sb00100000, 8'sb00100001, 8'sb00011110, 8'sb00101011, 8'sb00101000, 8'sb00111110, 8'sb00100100, 8'sb00010101, 8'sb11110100, 8'sb00000110, 8'sb00000110, 8'sb00101010, 8'sb00000010, 8'sb11101110, 8'sb11111110, 8'sb11111111, 8'sb11111111, 8'sb00001110, 8'sb00011101, 8'sb00110010, 8'sb00100000, 8'sb11111011, 8'sb11101010, 8'sb00100100, 8'sb11111011, 8'sb00101010, 8'sb11101111, 8'sb11111011, 8'sb00011111, 8'sb00010011, 8'sb00000111, 8'sb11110110, 8'sb00000001, 8'sb00011010, 8'sb11111000, 8'sb11111010, 8'sb00000010, 8'sb00000111, 8'sb11111101, 8'sb00000000, 8'sb11000010, 8'sb11010000, 8'sb11011000, 8'sb11100100, 8'sb11010001, 8'sb11011101, 8'sb11101100, 8'sb11100000, 8'sb11011111, 8'sb11110011, 8'sb11110000, 8'sb11111100,
    8'sb11111011, 8'sb11111101, 8'sb00001000, 8'sb00100010, 8'sb00100101, 8'sb00011110, 8'sb11111010, 8'sb00011000, 8'sb00000111, 8'sb01000000, 8'sb01000001, 8'sb00010101, 8'sb00000100, 8'sb11111101, 8'sb00001010, 8'sb00010100, 8'sb00101010, 8'sb00110000, 8'sb00010111, 8'sb11110011, 8'sb11111101, 8'sb00001100, 8'sb00010111, 8'sb00001100, 8'sb00001100, 8'sb00010111, 8'sb00000011, 8'sb11110101, 8'sb00001100, 8'sb00001000, 8'sb00011110, 8'sb00001110, 8'sb00000010, 8'sb11011100, 8'sb11101110, 8'sb00000011, 8'sb11100011, 8'sb11101110, 8'sb11111001, 8'sb00000111, 8'sb11110100, 8'sb11101001, 8'sb00010010, 8'sb00011111, 8'sb00001000, 8'sb00010001, 8'sb11111111, 8'sb11111110, 8'sb11110001, 8'sb11100100, 8'sb11100001, 8'sb11100000, 8'sb11100001, 8'sb11110110, 8'sb11111011, 8'sb00001110, 8'sb00101010, 8'sb00001010, 8'sb00011011, 8'sb00000011, 8'sb00001011, 8'sb11100111, 8'sb11101001, 8'sb11111010, 8'sb00000100, 8'sb11111000, 8'sb11111001, 8'sb11100101, 8'sb11100011, 8'sb11111100, 8'sb01000001, 8'sb00100001, 8'sb00010001, 8'sb00010011, 8'sb11111111, 8'sb11110001, 8'sb00010011, 8'sb01000100, 8'sb00101111, 8'sb00010100, 8'sb00011110, 8'sb00011011, 8'sb00001100, 8'sb11110101, 8'sb00110101, 8'sb00101010, 8'sb00001011, 8'sb00000001, 8'sb00000011, 8'sb00000010, 8'sb11110100, 8'sb00010010, 8'sb00010001, 8'sb00001100, 8'sb00001010, 8'sb00010001, 8'sb00010011, 8'sb11110110, 8'sb00011101, 8'sb00011111, 8'sb00001010, 8'sb00001101, 8'sb00001000, 8'sb00000001, 8'sb11100100, 8'sb00010111, 8'sb11111001, 8'sb00010101, 8'sb00011000, 8'sb00100000, 8'sb11101101, 8'sb10111110, 8'sb11110010, 8'sb11101101, 8'sb11111101, 8'sb00000101, 8'sb11110010, 8'sb11101001, 8'sb00010001, 8'sb00100110, 8'sb11110000, 8'sb00001110, 8'sb00010011, 8'sb00000001, 8'sb11101011, 8'sb11101110, 8'sb00011010, 8'sb11111110, 8'sb11101000, 8'sb11110000, 8'sb11111101, 8'sb00000000, 8'sb00101100, 8'sb00010111, 8'sb11111010, 8'sb11110011, 8'sb11101101, 8'sb11010001, 8'sb11100001, 8'sb00011110, 8'sb00000010, 8'sb10101111, 8'sb11011000, 8'sb11101101, 8'sb00000001, 8'sb00001111, 8'sb00010010, 8'sb00010011, 8'sb11110010, 8'sb11011001, 8'sb10111100, 8'sb10011001, 8'sb11000011, 8'sb00010111, 8'sb00001000, 8'sb11000010, 8'sb00010100, 8'sb00001110, 8'sb11111100, 8'sb11111000, 8'sb11110111, 8'sb00000010, 8'sb11110001, 8'sb11011001, 8'sb11001000, 8'sb10110010, 8'sb11101101, 8'sb00011111, 8'sb00000100, 8'sb11111101, 8'sb00011011, 8'sb00010001, 8'sb11110110, 8'sb11101101, 8'sb11101011, 8'sb11110001, 8'sb11100110, 8'sb11011111, 8'sb11100101, 8'sb11011100, 8'sb11111000, 8'sb00011111, 8'sb11110100, 8'sb11110110, 8'sb11010001, 8'sb00000001, 8'sb00001001, 8'sb00000111, 8'sb11111011, 8'sb11101010, 8'sb11100100, 8'sb11111010, 8'sb00000110, 8'sb00001001, 8'sb00000110, 8'sb00000111,
    8'sb11111011, 8'sb11110111, 8'sb11111111, 8'sb00011001, 8'sb00101110, 8'sb00101111, 8'sb00101001, 8'sb11110100, 8'sb00110110, 8'sb00110011, 8'sb00110001, 8'sb00011001, 8'sb00000101, 8'sb00000110, 8'sb00000000, 8'sb00100111, 8'sb00001101, 8'sb00001100, 8'sb00110010, 8'sb00110110, 8'sb00110110, 8'sb00100011, 8'sb00011001, 8'sb00011011, 8'sb00001110, 8'sb00101100, 8'sb00011100, 8'sb00011010, 8'sb11111101, 8'sb00000101, 8'sb11100100, 8'sb11101110, 8'sb11110110, 8'sb00001001, 8'sb11111101, 8'sb00000010, 8'sb00010111, 8'sb00011010, 8'sb00011100, 8'sb00011000, 8'sb00000111, 8'sb00100010, 8'sb00000101, 8'sb11101110, 8'sb00000000, 8'sb11111101, 8'sb11101100, 8'sb11110001, 8'sb11110100, 8'sb11111000, 8'sb11011111, 8'sb11110010, 8'sb11100111, 8'sb11111001, 8'sb00011000, 8'sb00010111, 8'sb00000001, 8'sb00000111, 8'sb11101100, 8'sb11111100, 8'sb11111011, 8'sb00001110, 8'sb00001011, 8'sb11101111, 8'sb11111011, 8'sb11111000, 8'sb11101111, 8'sb11011001, 8'sb00011000, 8'sb11110110, 8'sb00001010, 8'sb11110110, 8'sb00000000, 8'sb00010011, 8'sb11111010, 8'sb11110000, 8'sb11111011, 8'sb11110000, 8'sb11111010, 8'sb11111010, 8'sb11110001, 8'sb11101010, 8'sb00110001, 8'sb00000101, 8'sb11111011, 8'sb11111010, 8'sb11110011, 8'sb00011010, 8'sb11111101, 8'sb11110111, 8'sb00010010, 8'sb11011100, 8'sb11101010, 8'sb11111011, 8'sb11111000, 8'sb00010000, 8'sb00110011, 8'sb11110111, 8'sb00000111, 8'sb00001011, 8'sb00001011, 8'sb00010101, 8'sb00011001, 8'sb00011100, 8'sb00011110, 8'sb11110110, 8'sb11111001, 8'sb11110111, 8'sb11111111, 8'sb00001111, 8'sb01000001, 8'sb00001110, 8'sb11011000, 8'sb00011001, 8'sb00001011, 8'sb00000010, 8'sb00001100, 8'sb00011111, 8'sb00010101, 8'sb00000110, 8'sb00010000, 8'sb11111100, 8'sb00000010, 8'sb00011111, 8'sb00110011, 8'sb00000100, 8'sb11011111, 8'sb00001010, 8'sb00011000, 8'sb00100010, 8'sb00010111, 8'sb00101110, 8'sb00010111, 8'sb00010011, 8'sb00010111, 8'sb00000001, 8'sb00001100, 8'sb00101110, 8'sb00011100, 8'sb11010110, 8'sb00001100, 8'sb00110000, 8'sb00011101, 8'sb00010010, 8'sb00101000, 8'sb00101000, 8'sb00101011, 8'sb00010101, 8'sb00001011, 8'sb00010001, 8'sb00001011, 8'sb00110001, 8'sb11111000, 8'sb00011001, 8'sb00000000, 8'sb01000000, 8'sb00001010, 8'sb11110100, 8'sb00010010, 8'sb00010110, 8'sb00000010, 8'sb00001101, 8'sb00000001, 8'sb00000011, 8'sb00001001, 8'sb00011101, 8'sb00000001, 8'sb00011100, 8'sb11111010, 8'sb00000000, 8'sb11010001, 8'sb11001010, 8'sb11000000, 8'sb11010111, 8'sb11100100, 8'sb11011001, 8'sb11100000, 8'sb11110101, 8'sb11111010, 8'sb00010010, 8'sb00010110, 8'sb11110010, 8'sb11110111, 8'sb11110101, 8'sb00000000, 8'sb11010110, 8'sb10110010, 8'sb11101001, 8'sb11111011, 8'sb11011111, 8'sb11110100, 8'sb11101101, 8'sb11011011, 8'sb11101100, 8'sb11110100, 8'sb11111000,
    8'sb11111101, 8'sb11111010, 8'sb11111100, 8'sb11110110, 8'sb00011011, 8'sb00010101, 8'sb00001101, 8'sb00100000, 8'sb11111111, 8'sb11110111, 8'sb11110011, 8'sb11110110, 8'sb00001000, 8'sb00001001, 8'sb11111010, 8'sb11110011, 8'sb00001011, 8'sb11111010, 8'sb11110111, 8'sb11111001, 8'sb00011100, 8'sb00011110, 8'sb00100010, 8'sb00010010, 8'sb00011010, 8'sb00010100, 8'sb00010101, 8'sb00001000, 8'sb11111000, 8'sb11110011, 8'sb11101001, 8'sb11111011, 8'sb00010101, 8'sb00100110, 8'sb00001011, 8'sb00010000, 8'sb00000111, 8'sb00000011, 8'sb00010010, 8'sb00100110, 8'sb00111111, 8'sb00010011, 8'sb00010011, 8'sb00000000, 8'sb00000110, 8'sb00010001, 8'sb00010010, 8'sb00011010, 8'sb11111101, 8'sb11100010, 8'sb11110111, 8'sb00000100, 8'sb00000010, 8'sb11111110, 8'sb00100111, 8'sb11111111, 8'sb00011010, 8'sb11111111, 8'sb00010000, 8'sb00100100, 8'sb00100001, 8'sb00101000, 8'sb11100100, 8'sb11011100, 8'sb11111111, 8'sb00000101, 8'sb11111011, 8'sb11101011, 8'sb00010100, 8'sb11101110, 8'sb00111110, 8'sb00001110, 8'sb00000000, 8'sb00010111, 8'sb00111000, 8'sb00110010, 8'sb10111110, 8'sb11100010, 8'sb00011010, 8'sb11110110, 8'sb11110110, 8'sb11101110, 8'sb11110000, 8'sb11100101, 8'sb01000001, 8'sb00010110, 8'sb00100001, 8'sb00101100, 8'sb00100110, 8'sb00010011, 8'sb10101011, 8'sb11100010, 8'sb00010010, 8'sb00000000, 8'sb00000011, 8'sb00010010, 8'sb11110100, 8'sb11011011, 8'sb00101011, 8'sb00001100, 8'sb00100100, 8'sb00101100, 8'sb00110100, 8'sb00000111, 8'sb11011101, 8'sb11000111, 8'sb00000101, 8'sb00001000, 8'sb11111110, 8'sb00101000, 8'sb00000100, 8'sb11011100, 8'sb00000011, 8'sb11100011, 8'sb11111100, 8'sb00010101, 8'sb00101011, 8'sb00001001, 8'sb11010111, 8'sb11011010, 8'sb11111111, 8'sb00000000, 8'sb00001101, 8'sb00011000, 8'sb00000010, 8'sb11010111, 8'sb00010011, 8'sb00010000, 8'sb11110101, 8'sb11110110, 8'sb00001010, 8'sb00001010, 8'sb11011010, 8'sb11111001, 8'sb00001100, 8'sb00100000, 8'sb00011111, 8'sb00010010, 8'sb00000000, 8'sb11001100, 8'sb11101100, 8'sb11101010, 8'sb11111110, 8'sb11101101, 8'sb11110111, 8'sb11110000, 8'sb11110010, 8'sb00001000, 8'sb00101111, 8'sb00011111, 8'sb00011111, 8'sb11111110, 8'sb00001000, 8'sb11100111, 8'sb00000110, 8'sb11011001, 8'sb00000001, 8'sb11101100, 8'sb11000010, 8'sb11011001, 8'sb11101111, 8'sb00100011, 8'sb00101011, 8'sb00100111, 8'sb00011000, 8'sb00000000, 8'sb00000111, 8'sb00011100, 8'sb11111010, 8'sb00011011, 8'sb00000110, 8'sb11101010, 8'sb11011111, 8'sb11110011, 8'sb00001000, 8'sb00000011, 8'sb00001101, 8'sb00001010, 8'sb11111111, 8'sb00000100, 8'sb11011100, 8'sb11111000, 8'sb00001001, 8'sb00000011, 8'sb00000110, 8'sb00000101, 8'sb00100001, 8'sb00000111, 8'sb00001110, 8'sb00000101, 8'sb00100001, 8'sb00101100, 8'sb00101010, 8'sb00010100, 8'sb11110100, 8'sb00000101,
    8'sb00000011, 8'sb11111011, 8'sb00001001, 8'sb00000010, 8'sb00000000, 8'sb00000100, 8'sb11110101, 8'sb00010000, 8'sb00010110, 8'sb00101011, 8'sb00001010, 8'sb00001011, 8'sb11111101, 8'sb00000001, 8'sb00001100, 8'sb00001100, 8'sb00011011, 8'sb00011110, 8'sb00010011, 8'sb00100100, 8'sb00101110, 8'sb00101010, 8'sb00100001, 8'sb00100111, 8'sb00011011, 8'sb11110001, 8'sb00000010, 8'sb00001000, 8'sb00001100, 8'sb00010001, 8'sb00001001, 8'sb00000100, 8'sb00011011, 8'sb00010000, 8'sb00000100, 8'sb00001100, 8'sb00001110, 8'sb00010111, 8'sb00010110, 8'sb00011111, 8'sb00100010, 8'sb00010101, 8'sb00011101, 8'sb11111101, 8'sb00001111, 8'sb00010000, 8'sb00010101, 8'sb00010001, 8'sb00001100, 8'sb00010111, 8'sb00010100, 8'sb00001000, 8'sb00011000, 8'sb00010011, 8'sb00010100, 8'sb00000111, 8'sb00001100, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00100100, 8'sb00011100, 8'sb00001001, 8'sb00000110, 8'sb11111101, 8'sb00010100, 8'sb00000001, 8'sb00011101, 8'sb11110011, 8'sb00111011, 8'sb00001010, 8'sb00000101, 8'sb11111110, 8'sb00001011, 8'sb00011001, 8'sb00001110, 8'sb11110100, 8'sb11101111, 8'sb11100111, 8'sb11111001, 8'sb00001001, 8'sb00110000, 8'sb11110101, 8'sb00010100, 8'sb11111111, 8'sb11101000, 8'sb11110100, 8'sb11101101, 8'sb00001100, 8'sb00001100, 8'sb11111110, 8'sb11111010, 8'sb11100001, 8'sb11000111, 8'sb10110110, 8'sb11111010, 8'sb00010000, 8'sb11110110, 8'sb11101100, 8'sb11100010, 8'sb11100011, 8'sb11100111, 8'sb00010010, 8'sb00000111, 8'sb11110101, 8'sb11111100, 8'sb00001110, 8'sb00001001, 8'sb11110011, 8'sb10111101, 8'sb00100011, 8'sb00010110, 8'sb11111110, 8'sb11011100, 8'sb11001001, 8'sb00000011, 8'sb00010000, 8'sb11011000, 8'sb11011100, 8'sb00001110, 8'sb00000111, 8'sb00001111, 8'sb11111000, 8'sb11000110, 8'sb00110000, 8'sb00100111, 8'sb00010010, 8'sb11110100, 8'sb11100000, 8'sb11101101, 8'sb11100101, 8'sb11100000, 8'sb00000100, 8'sb00001001, 8'sb00010000, 8'sb00001011, 8'sb11011001, 8'sb10110100, 8'sb00010011, 8'sb00001100, 8'sb11111010, 8'sb00001010, 8'sb00000011, 8'sb00001110, 8'sb00010110, 8'sb00011011, 8'sb00001011, 8'sb00100101, 8'sb00011011, 8'sb00010100, 8'sb11000001, 8'sb11100010, 8'sb00000111, 8'sb00101011, 8'sb00001110, 8'sb00001001, 8'sb11110100, 8'sb00010000, 8'sb00010011, 8'sb00100000, 8'sb00100001, 8'sb00100001, 8'sb00000110, 8'sb11111110, 8'sb11010001, 8'sb11110010, 8'sb00000101, 8'sb00111100, 8'sb00000000, 8'sb00010101, 8'sb00100010, 8'sb00011111, 8'sb00111010, 8'sb00101000, 8'sb00011111, 8'sb00001000, 8'sb11111111, 8'sb00011001, 8'sb11111110, 8'sb11110011, 8'sb00001010, 8'sb11110111, 8'sb11101110, 8'sb11101101, 8'sb00001101, 8'sb00100001, 8'sb00100011, 8'sb00100010, 8'sb01001000, 8'sb00111100, 8'sb00101010, 8'sb00110000, 8'sb00001001, 8'sb11111101,
    8'sb11111011, 8'sb11110100, 8'sb00001100, 8'sb11111101, 8'sb11111101, 8'sb00001100, 8'sb00100010, 8'sb00000101, 8'sb11101011, 8'sb00011101, 8'sb00000001, 8'sb00000000, 8'sb00000100, 8'sb00000011, 8'sb00000100, 8'sb11101100, 8'sb00000011, 8'sb11111000, 8'sb11011001, 8'sb11101010, 8'sb00000101, 8'sb11111110, 8'sb11111111, 8'sb00001100, 8'sb11110001, 8'sb00001010, 8'sb11101111, 8'sb11110010, 8'sb00001011, 8'sb11110010, 8'sb11001100, 8'sb11010011, 8'sb11101011, 8'sb11100101, 8'sb00010100, 8'sb00000100, 8'sb00000010, 8'sb11101111, 8'sb11111111, 8'sb11111010, 8'sb00100011, 8'sb00010111, 8'sb11101110, 8'sb11011100, 8'sb11100111, 8'sb11110100, 8'sb11101010, 8'sb00001101, 8'sb00011010, 8'sb11110100, 8'sb11010101, 8'sb11110101, 8'sb11111010, 8'sb00001001, 8'sb00101011, 8'sb00011011, 8'sb11110001, 8'sb11010111, 8'sb11011100, 8'sb11100111, 8'sb11110010, 8'sb00011011, 8'sb00101100, 8'sb11011110, 8'sb11101010, 8'sb00001101, 8'sb00011000, 8'sb00010100, 8'sb00101000, 8'sb00100001, 8'sb00001111, 8'sb11011101, 8'sb11101100, 8'sb11101100, 8'sb11111011, 8'sb00001000, 8'sb00101100, 8'sb00000101, 8'sb11111001, 8'sb00000110, 8'sb00000000, 8'sb00010100, 8'sb00001111, 8'sb00010111, 8'sb11110000, 8'sb11101100, 8'sb11011111, 8'sb11111101, 8'sb11111010, 8'sb11110110, 8'sb00101101, 8'sb00001010, 8'sb11111001, 8'sb00000101, 8'sb00010110, 8'sb00100111, 8'sb00101011, 8'sb11010100, 8'sb00000111, 8'sb00010010, 8'sb11000001, 8'sb11100111, 8'sb11101000, 8'sb00001110, 8'sb00010110, 8'sb00001110, 8'sb11110100, 8'sb11111000, 8'sb11101011, 8'sb11101011, 8'sb11111001, 8'sb10111101, 8'sb11110000, 8'sb11101101, 8'sb11010001, 8'sb11011100, 8'sb00010011, 8'sb00100110, 8'sb00100010, 8'sb11101010, 8'sb11110001, 8'sb11110011, 8'sb11111001, 8'sb11110011, 8'sb11110110, 8'sb11010100, 8'sb11101101, 8'sb11011110, 8'sb11000110, 8'sb11101111, 8'sb00100010, 8'sb00101010, 8'sb00001110, 8'sb11001110, 8'sb11101110, 8'sb11110010, 8'sb11111011, 8'sb00000101, 8'sb11111000, 8'sb00001001, 8'sb11111110, 8'sb11010011, 8'sb11010010, 8'sb00000011, 8'sb00010010, 8'sb00010111, 8'sb11110010, 8'sb11111000, 8'sb11011101, 8'sb11101110, 8'sb00000001, 8'sb00000010, 8'sb11000111, 8'sb11101100, 8'sb00001110, 8'sb11101001, 8'sb11011110, 8'sb11110101, 8'sb00001010, 8'sb00001111, 8'sb00010001, 8'sb00001000, 8'sb11111101, 8'sb11110001, 8'sb11101001, 8'sb11011010, 8'sb11110011, 8'sb11111010, 8'sb11110110, 8'sb11011001, 8'sb11101101, 8'sb11011101, 8'sb11111010, 8'sb00011010, 8'sb00010011, 8'sb00001001, 8'sb11110010, 8'sb11100110, 8'sb11110011, 8'sb11101001, 8'sb11111001, 8'sb00000001, 8'sb11111001, 8'sb11110100, 8'sb11011100, 8'sb11010011, 8'sb11010100, 8'sb11010101, 8'sb11010111, 8'sb10101110, 8'sb11000111, 8'sb11000001, 8'sb11000100, 8'sb00011001, 8'sb00001101, 8'sb00001010,
    8'sb00000010, 8'sb11111011, 8'sb00000011, 8'sb11100111, 8'sb11011111, 8'sb11010010, 8'sb11001110, 8'sb11110111, 8'sb11011000, 8'sb10111101, 8'sb11001011, 8'sb11101001, 8'sb00000100, 8'sb00000110, 8'sb11111011, 8'sb11100001, 8'sb11011110, 8'sb11001001, 8'sb11000001, 8'sb11001000, 8'sb10010001, 8'sb10111111, 8'sb11100001, 8'sb00000000, 8'sb11100100, 8'sb11100010, 8'sb11101011, 8'sb11111110, 8'sb00001010, 8'sb00000000, 8'sb11100100, 8'sb11010110, 8'sb11000100, 8'sb10011100, 8'sb10100000, 8'sb11000000, 8'sb11011100, 8'sb11101111, 8'sb11101100, 8'sb11110110, 8'sb00001000, 8'sb11101011, 8'sb00010000, 8'sb00111011, 8'sb11110110, 8'sb00000101, 8'sb00011100, 8'sb11111001, 8'sb11111010, 8'sb11111000, 8'sb00000010, 8'sb00000000, 8'sb00001010, 8'sb11110101, 8'sb11101111, 8'sb00001010, 8'sb00011001, 8'sb00000111, 8'sb00001011, 8'sb00001110, 8'sb00011011, 8'sb00111000, 8'sb00111011, 8'sb00011000, 8'sb11111001, 8'sb11111101, 8'sb00000011, 8'sb00000101, 8'sb11100100, 8'sb00001111, 8'sb11110101, 8'sb00100011, 8'sb11110010, 8'sb00011001, 8'sb00101001, 8'sb00011001, 8'sb00001000, 8'sb00001111, 8'sb00000110, 8'sb00001010, 8'sb00000101, 8'sb11100001, 8'sb11010101, 8'sb00001110, 8'sb00110001, 8'sb00001001, 8'sb11110000, 8'sb00001100, 8'sb11111011, 8'sb11110110, 8'sb11111000, 8'sb00001101, 8'sb00010101, 8'sb00001100, 8'sb00010001, 8'sb11100100, 8'sb11110111, 8'sb01001001, 8'sb00001000, 8'sb00010011, 8'sb00000011, 8'sb00010111, 8'sb00001010, 8'sb00001101, 8'sb00011100, 8'sb00010010, 8'sb00011110, 8'sb00100100, 8'sb00010001, 8'sb00000110, 8'sb00000010, 8'sb01001111, 8'sb00010000, 8'sb00011011, 8'sb00001001, 8'sb00000111, 8'sb00011010, 8'sb00010110, 8'sb00011000, 8'sb00000111, 8'sb00011111, 8'sb00010101, 8'sb00001110, 8'sb00001100, 8'sb11101101, 8'sb00111010, 8'sb11111111, 8'sb00101011, 8'sb00000010, 8'sb11100011, 8'sb11010101, 8'sb11011100, 8'sb11011011, 8'sb11110000, 8'sb11111011, 8'sb11111101, 8'sb00000010, 8'sb00001111, 8'sb11111111, 8'sb00101011, 8'sb11110110, 8'sb00011001, 8'sb11101001, 8'sb11010110, 8'sb11011010, 8'sb11010110, 8'sb11100011, 8'sb11011111, 8'sb11100111, 8'sb11011111, 8'sb11101011, 8'sb11101001, 8'sb00000110, 8'sb11110011, 8'sb00000011, 8'sb00010100, 8'sb11110011, 8'sb11110011, 8'sb11110010, 8'sb00000000, 8'sb11101011, 8'sb11011100, 8'sb11100010, 8'sb11011001, 8'sb11011010, 8'sb11100010, 8'sb11111000, 8'sb11110000, 8'sb00001001, 8'sb00000111, 8'sb00111010, 8'sb00100111, 8'sb00000011, 8'sb00000110, 8'sb00000000, 8'sb11110111, 8'sb00010101, 8'sb11111011, 8'sb00001010, 8'sb00010000, 8'sb00001111, 8'sb00011101, 8'sb11111001, 8'sb11111001, 8'sb11111100, 8'sb00100001, 8'sb00101011, 8'sb00101110, 8'sb00111001, 8'sb00111010, 8'sb00110011, 8'sb00101001, 8'sb00101011, 8'sb00010001, 8'sb00000000, 8'sb11111111,
    8'sb00000110, 8'sb11111011, 8'sb11111100, 8'sb11111100, 8'sb00001011, 8'sb00010110, 8'sb00001100, 8'sb00001011, 8'sb00001101, 8'sb00010000, 8'sb00000010, 8'sb00001101, 8'sb11111111, 8'sb00000101, 8'sb11110111, 8'sb11111001, 8'sb11011011, 8'sb11100101, 8'sb11111011, 8'sb11110100, 8'sb00010100, 8'sb00101000, 8'sb00011001, 8'sb00000001, 8'sb11111101, 8'sb11100110, 8'sb00010011, 8'sb00011101, 8'sb00000110, 8'sb00000011, 8'sb11101000, 8'sb11101110, 8'sb11111111, 8'sb11110000, 8'sb11111111, 8'sb00000100, 8'sb11111111, 8'sb00000101, 8'sb11111011, 8'sb00000110, 8'sb11110110, 8'sb00101011, 8'sb11101001, 8'sb00100001, 8'sb00010011, 8'sb00001111, 8'sb00000100, 8'sb00001011, 8'sb00010110, 8'sb00011110, 8'sb00010010, 8'sb00010001, 8'sb00011010, 8'sb00000101, 8'sb00000101, 8'sb00001000, 8'sb00101111, 8'sb00000010, 8'sb00001011, 8'sb00000101, 8'sb00011001, 8'sb00001111, 8'sb00100111, 8'sb00101111, 8'sb00011100, 8'sb00000001, 8'sb11111000, 8'sb00000110, 8'sb11110101, 8'sb11100110, 8'sb00111001, 8'sb00100101, 8'sb00010001, 8'sb00011001, 8'sb00010011, 8'sb00011111, 8'sb00010111, 8'sb11110000, 8'sb11110010, 8'sb00000111, 8'sb11111010, 8'sb11111100, 8'sb11110000, 8'sb11110010, 8'sb00100110, 8'sb00001111, 8'sb11110010, 8'sb00001111, 8'sb11111101, 8'sb00000100, 8'sb11001101, 8'sb11001100, 8'sb11110001, 8'sb11111010, 8'sb00000100, 8'sb00011001, 8'sb00001111, 8'sb11101011, 8'sb00001000, 8'sb11110011, 8'sb11111110, 8'sb11111000, 8'sb11101001, 8'sb11011011, 8'sb11010110, 8'sb11010111, 8'sb11011100, 8'sb11110010, 8'sb00001110, 8'sb00011101, 8'sb00101010, 8'sb11111101, 8'sb11110111, 8'sb11100001, 8'sb00010010, 8'sb11110111, 8'sb11011100, 8'sb11100110, 8'sb10110001, 8'sb11010001, 8'sb11111000, 8'sb00000100, 8'sb00001100, 8'sb00000110, 8'sb11110101, 8'sb11111111, 8'sb00011011, 8'sb11100100, 8'sb11101100, 8'sb11101110, 8'sb11100010, 8'sb11011110, 8'sb10111011, 8'sb00001001, 8'sb00010101, 8'sb00001110, 8'sb00001101, 8'sb11111101, 8'sb11110011, 8'sb11110011, 8'sb11111111, 8'sb11110101, 8'sb00001001, 8'sb00001100, 8'sb00000001, 8'sb00000111, 8'sb00101010, 8'sb00100111, 8'sb00001110, 8'sb11110100, 8'sb11110110, 8'sb11111001, 8'sb00101010, 8'sb00001101, 8'sb11111000, 8'sb11010000, 8'sb11111110, 8'sb11110111, 8'sb00011011, 8'sb00100011, 8'sb00011010, 8'sb00100110, 8'sb00010110, 8'sb11101110, 8'sb11111010, 8'sb00000001, 8'sb11110110, 8'sb11101111, 8'sb11110111, 8'sb00000011, 8'sb11110101, 8'sb00000100, 8'sb00011101, 8'sb11111100, 8'sb00000001, 8'sb00000111, 8'sb00011001, 8'sb11111010, 8'sb00001010, 8'sb11111000, 8'sb00000010, 8'sb11111110, 8'sb00001011, 8'sb11111100, 8'sb00000010, 8'sb00010011, 8'sb01011001, 8'sb00110110, 8'sb00101110, 8'sb01010011, 8'sb01010100, 8'sb01011111, 8'sb01000011, 8'sb00111010, 8'sb00001010, 8'sb00000011,
    8'sb00001001, 8'sb00000100, 8'sb00000101, 8'sb11110010, 8'sb11011111, 8'sb11101000, 8'sb11011110, 8'sb00011001, 8'sb00010001, 8'sb11010000, 8'sb11010110, 8'sb11101011, 8'sb00001100, 8'sb00001100, 8'sb11111101, 8'sb00001001, 8'sb11111010, 8'sb11111101, 8'sb00001101, 8'sb00001101, 8'sb00000110, 8'sb00000000, 8'sb11111000, 8'sb11100100, 8'sb11001010, 8'sb11011101, 8'sb11110001, 8'sb11110001, 8'sb11111111, 8'sb00000111, 8'sb00011000, 8'sb00100011, 8'sb00000101, 8'sb00011011, 8'sb00010110, 8'sb00000111, 8'sb11110110, 8'sb11100101, 8'sb11101000, 8'sb11010010, 8'sb11101010, 8'sb00010011, 8'sb00010110, 8'sb00110001, 8'sb00001000, 8'sb00001011, 8'sb00001011, 8'sb00001110, 8'sb00000100, 8'sb00011000, 8'sb00011100, 8'sb00001001, 8'sb11101110, 8'sb11011111, 8'sb11100000, 8'sb11110100, 8'sb11100100, 8'sb00001111, 8'sb00010101, 8'sb00010100, 8'sb00001010, 8'sb11111000, 8'sb00000011, 8'sb00011110, 8'sb00011100, 8'sb00010111, 8'sb00011011, 8'sb11111001, 8'sb11011110, 8'sb11111011, 8'sb11101101, 8'sb00110010, 8'sb00010110, 8'sb00001111, 8'sb00000100, 8'sb11101011, 8'sb00001001, 8'sb00100111, 8'sb00001111, 8'sb00011100, 8'sb00110011, 8'sb00100011, 8'sb11011011, 8'sb00010100, 8'sb00000010, 8'sb00100101, 8'sb00010000, 8'sb11110010, 8'sb11101110, 8'sb11101101, 8'sb00000011, 8'sb00110000, 8'sb00100011, 8'sb00011100, 8'sb00100110, 8'sb00000100, 8'sb11101001, 8'sb00010110, 8'sb11111100, 8'sb00001010, 8'sb11110011, 8'sb11101010, 8'sb11101000, 8'sb11101100, 8'sb00001010, 8'sb00100000, 8'sb00000100, 8'sb00011010, 8'sb11111110, 8'sb11100001, 8'sb11011110, 8'sb00001111, 8'sb00011010, 8'sb00010001, 8'sb11111100, 8'sb11101110, 8'sb11111101, 8'sb00001010, 8'sb00011011, 8'sb00000110, 8'sb00000101, 8'sb11101010, 8'sb11100011, 8'sb11110110, 8'sb11011110, 8'sb00000100, 8'sb00011110, 8'sb11111100, 8'sb11101110, 8'sb11110110, 8'sb00001011, 8'sb00001101, 8'sb00000101, 8'sb11110010, 8'sb11111100, 8'sb11110111, 8'sb11111011, 8'sb00001110, 8'sb11110100, 8'sb00100001, 8'sb11110101, 8'sb11110010, 8'sb00000001, 8'sb00000111, 8'sb11110011, 8'sb11101010, 8'sb11110111, 8'sb00000010, 8'sb11111111, 8'sb00000111, 8'sb00000010, 8'sb11111000, 8'sb00000101, 8'sb11101110, 8'sb00001010, 8'sb00011000, 8'sb11111111, 8'sb00001110, 8'sb11111100, 8'sb00000000, 8'sb11110110, 8'sb00000100, 8'sb11111000, 8'sb00000000, 8'sb00001001, 8'sb00010101, 8'sb00000100, 8'sb11100011, 8'sb11110100, 8'sb00001110, 8'sb00100100, 8'sb00011011, 8'sb00000100, 8'sb00010110, 8'sb00010100, 8'sb00000010, 8'sb00011001, 8'sb00010010, 8'sb00010101, 8'sb00000001, 8'sb11111010, 8'sb00000100, 8'sb00000111, 8'sb00000111, 8'sb00011101, 8'sb01010000, 8'sb01011111, 8'sb01001101, 8'sb01010001, 8'sb01010001, 8'sb01000101, 8'sb00111000, 8'sb00110110, 8'sb00010111, 8'sb00011101, 8'sb11110111,
    8'sb11111011, 8'sb11110100, 8'sb11110110, 8'sb11010010, 8'sb11101010, 8'sb00001001, 8'sb11101101, 8'sb11101011, 8'sb00000101, 8'sb11001011, 8'sb11000111, 8'sb11101000, 8'sb00000111, 8'sb11110110, 8'sb00001010, 8'sb11110100, 8'sb00000010, 8'sb00011000, 8'sb00100000, 8'sb01001100, 8'sb00010011, 8'sb00010011, 8'sb00000110, 8'sb11111001, 8'sb00001000, 8'sb11010111, 8'sb00010010, 8'sb00000101, 8'sb11111110, 8'sb00001010, 8'sb00100100, 8'sb00101111, 8'sb00100110, 8'sb00011000, 8'sb00001010, 8'sb00000010, 8'sb00000011, 8'sb00000001, 8'sb11111001, 8'sb00000111, 8'sb11101000, 8'sb11100010, 8'sb00011111, 8'sb00110010, 8'sb01000010, 8'sb00011100, 8'sb00000001, 8'sb00001010, 8'sb00100101, 8'sb00001001, 8'sb11101011, 8'sb11101001, 8'sb11110111, 8'sb00000101, 8'sb11010110, 8'sb11111100, 8'sb00101010, 8'sb00110100, 8'sb00010010, 8'sb11100011, 8'sb11001010, 8'sb11011001, 8'sb00000001, 8'sb00011001, 8'sb00000111, 8'sb00001000, 8'sb00000000, 8'sb11110001, 8'sb11101111, 8'sb11011011, 8'sb00100111, 8'sb00100101, 8'sb10111100, 8'sb10110100, 8'sb10110101, 8'sb11011010, 8'sb00010010, 8'sb11111000, 8'sb00010000, 8'sb00000110, 8'sb00000110, 8'sb11101011, 8'sb11010010, 8'sb11000010, 8'sb00011010, 8'sb11100100, 8'sb11000011, 8'sb11100100, 8'sb00000001, 8'sb00100110, 8'sb00010110, 8'sb11011001, 8'sb11100111, 8'sb11110010, 8'sb11010111, 8'sb11101100, 8'sb00000001, 8'sb11110111, 8'sb00100111, 8'sb00010010, 8'sb00001010, 8'sb00010000, 8'sb00011011, 8'sb00011101, 8'sb11111000, 8'sb11100010, 8'sb11101110, 8'sb00000011, 8'sb00000100, 8'sb00100011, 8'sb00101111, 8'sb01010100, 8'sb00100001, 8'sb01001100, 8'sb00110001, 8'sb11110110, 8'sb00000011, 8'sb11111101, 8'sb11110111, 8'sb11110001, 8'sb00011110, 8'sb00100101, 8'sb00110010, 8'sb00100100, 8'sb00001000, 8'sb00111000, 8'sb00000110, 8'sb00111011, 8'sb00011010, 8'sb00000001, 8'sb00000111, 8'sb00010111, 8'sb00010110, 8'sb00001101, 8'sb00010000, 8'sb00000010, 8'sb00001100, 8'sb00000110, 8'sb11110001, 8'sb00010000, 8'sb00010010, 8'sb00111011, 8'sb00001010, 8'sb11101111, 8'sb00000110, 8'sb00010011, 8'sb00011000, 8'sb00001000, 8'sb00000011, 8'sb00000011, 8'sb11111101, 8'sb11111011, 8'sb11101001, 8'sb00010010, 8'sb11110110, 8'sb00111000, 8'sb11111101, 8'sb00000111, 8'sb00000001, 8'sb00010000, 8'sb11111111, 8'sb00000110, 8'sb00000000, 8'sb00001011, 8'sb11101101, 8'sb11101111, 8'sb11101100, 8'sb11110111, 8'sb00000101, 8'sb00110110, 8'sb00011010, 8'sb11111010, 8'sb00000000, 8'sb11111100, 8'sb11111101, 8'sb11111101, 8'sb11111011, 8'sb11101110, 8'sb11110000, 8'sb11111010, 8'sb00000011, 8'sb11101111, 8'sb00001001, 8'sb11100110, 8'sb11100110, 8'sb11011111, 8'sb11100101, 8'sb11101001, 8'sb11101110, 8'sb11110011, 8'sb00011001, 8'sb00001010, 8'sb11101110, 8'sb11110000, 8'sb11110110, 8'sb11111101,
    8'sb11111110, 8'sb00000001, 8'sb11110000, 8'sb11110011, 8'sb11101011, 8'sb11100010, 8'sb11010100, 8'sb00011111, 8'sb00100000, 8'sb11000110, 8'sb11010101, 8'sb11101110, 8'sb11111011, 8'sb11111000, 8'sb00000011, 8'sb00100000, 8'sb00010010, 8'sb11111010, 8'sb00100010, 8'sb00000001, 8'sb00000101, 8'sb11110011, 8'sb00000110, 8'sb11110010, 8'sb11100100, 8'sb11011011, 8'sb11110000, 8'sb00000011, 8'sb00000001, 8'sb00011000, 8'sb00111001, 8'sb00010011, 8'sb00000101, 8'sb00010000, 8'sb00001000, 8'sb11111111, 8'sb00000110, 8'sb11111010, 8'sb00000111, 8'sb00010011, 8'sb11111100, 8'sb11101000, 8'sb00101111, 8'sb00000100, 8'sb11111010, 8'sb00001000, 8'sb00010000, 8'sb00101111, 8'sb00010010, 8'sb00001000, 8'sb00010101, 8'sb00011010, 8'sb00001111, 8'sb00001000, 8'sb00000000, 8'sb00001011, 8'sb00100111, 8'sb00000111, 8'sb11111100, 8'sb00001100, 8'sb00010101, 8'sb00100001, 8'sb00010101, 8'sb00010000, 8'sb00000100, 8'sb00000110, 8'sb11110101, 8'sb00000011, 8'sb11011111, 8'sb00010011, 8'sb11111010, 8'sb11010011, 8'sb11100000, 8'sb11101100, 8'sb11011111, 8'sb11001010, 8'sb10110110, 8'sb11110110, 8'sb11100011, 8'sb11001000, 8'sb11000000, 8'sb11001100, 8'sb11110001, 8'sb00011010, 8'sb00011000, 8'sb11010101, 8'sb10010001, 8'sb10001000, 8'sb10010010, 8'sb10100101, 8'sb11011100, 8'sb00001001, 8'sb11101101, 8'sb11110110, 8'sb11100101, 8'sb11001111, 8'sb11111101, 8'sb00110100, 8'sb11011111, 8'sb11101101, 8'sb11100100, 8'sb11100010, 8'sb11111010, 8'sb11111111, 8'sb00111000, 8'sb00100110, 8'sb00001001, 8'sb00011010, 8'sb00010001, 8'sb00001110, 8'sb00001100, 8'sb00110001, 8'sb11100100, 8'sb00000011, 8'sb00011000, 8'sb00011110, 8'sb00011100, 8'sb00010100, 8'sb00100100, 8'sb00010011, 8'sb00000101, 8'sb00000000, 8'sb00001011, 8'sb11111011, 8'sb00011101, 8'sb00110010, 8'sb11110110, 8'sb00010000, 8'sb00011001, 8'sb00011010, 8'sb00011110, 8'sb00001100, 8'sb00010011, 8'sb00000101, 8'sb00000111, 8'sb00001010, 8'sb00000101, 8'sb00000011, 8'sb01001110, 8'sb00101000, 8'sb11110101, 8'sb00001110, 8'sb00100100, 8'sb00010011, 8'sb00001101, 8'sb00001100, 8'sb00001111, 8'sb00010100, 8'sb00000100, 8'sb00000001, 8'sb00000111, 8'sb11111001, 8'sb00100001, 8'sb00011001, 8'sb00000011, 8'sb11011110, 8'sb00101110, 8'sb00001001, 8'sb11110001, 8'sb11111100, 8'sb00000011, 8'sb11110001, 8'sb11111100, 8'sb11100110, 8'sb11110100, 8'sb11111001, 8'sb00010110, 8'sb00100001, 8'sb00001001, 8'sb11100001, 8'sb00000111, 8'sb00000000, 8'sb00000101, 8'sb11110110, 8'sb00000010, 8'sb11111100, 8'sb11101001, 8'sb11100111, 8'sb11101010, 8'sb11100010, 8'sb00000000, 8'sb00011011, 8'sb00001001, 8'sb11110100, 8'sb11100110, 8'sb00000011, 8'sb00011011, 8'sb00011001, 8'sb11110110, 8'sb00001111, 8'sb11101111, 8'sb11110110, 8'sb11100000, 8'sb11110000, 8'sb00001101, 8'sb11110111
    };
    
    dense_layer #(
        .NEURON_NB(HL_neurons),
        .IN_SIZE(averaged_pixels_nr), 
        .WIDTH(WIDTH),
        .WIDTH_IN(WIDTH),
        .WIDTH_OUT(4*WIDTH)
    ) hidden_dense (
        .clk(clk), 
        .dense_go(hidden_go), 
        .reset(reset),
        .dense_in(hidden_in), 
        .weights(weights_HL_param), 
        .biases(biases_HL_param),
        .dense_out(dense_out), 
        .dense_done(dense_done)
    ); //Dense layer
    
    ReLU_layer #(
        .NEURON_NB(HL_neurons),
        .IN_SIZE(averaged_pixels_nr),
        .WIDTH(4*WIDTH)
    ) ReLU_hidden_layer (
        .clk(clk),
        .reset(reset),
        .relu_go(dense_done),
        .data_in_array(dense_out),
        .relu_layer_done(hidden_done),
        .data_out_array(hidden_out)
    );               

endmodule
