module hidden_layer_param (
    output reg signed [8*30*196-1:0] weights_HL, // Declare output as a flattened 1D array for weights
    output reg signed [8*30-1:0] biases_HL // Declare output as a flattened 1D array for biases
);

    // Local parameters for initialized weights and biases
    localparam signed [8*30*196-1:0] weights_HL_param = {
    8'sd11, 8'sd10, 8'sd11, 8'sd11, 8'sd12, 8'sd11, 8'sd14, 8'sd13, 8'sd11, 8'sd11, 8'sd13, 8'sd12, 8'sd14, 8'sd12, 8'sd10, 8'sd10, 8'sd11, 8'sd13, 8'sd16, 8'sd17, 8'sd21, 8'sd18, 8'sd17, 8'sd17, 8'sd16, 8'sd17, 8'sd13, 8'sd10, 8'sd11, 8'sd13, 8'sd12, 8'sd13, 8'sd9, 8'sd18, 8'sd23, 8'sd25, 8'sd23, 8'sd25, 8'sd20, 8'sd11, 8'sd13, 8'sd15, 8'sd14, 8'sd11, 8'sd13, 8'sd12, 8'sd13, 8'sd16, 8'sd17, 8'sd21, 8'sd8, 8'sd24, 8'sd19, 8'sd16, 8'sd22, 8'sd13, 8'sd13, 8'sd12, 8'sd14, 8'sd15, 8'sd15, 8'sd11, 8'sd9, 8'sd13, 8'sd22, 8'sd15, 8'sd24, 8'sd26, 8'sd35, 8'sd18, 8'sd12, 8'sd14, 8'sd15, 8'sd8, 8'sd6, 8'sd13, 8'sd8, 8'sd19, -8'sd8, -8'sd1, 8'sd11, 8'sd32, 8'sd36, 8'sd14, 8'sd14, 8'sd14, 8'sd13, 8'sd10, 8'sd10, 8'sd2, 8'sd28, 8'sd4, -8'sd10, -8'sd1, 8'sd3, 8'sd23, 8'sd19, 8'sd11, 8'sd11, 8'sd14, 8'sd4, 8'sd3, 8'sd8, 8'sd16, 8'sd27, 8'sd10, -8'sd8, -8'sd15, 8'sd7, 8'sd10, 8'sd14, 8'sd9, 8'sd13, 8'sd14, 8'sd0, -8'sd4, 8'sd10, 8'sd20, 8'sd26, -8'sd6, -8'sd10, -8'sd4, 8'sd8, 8'sd19, 8'sd12, 8'sd10, 8'sd12, 8'sd13, 8'sd12, 8'sd28, 8'sd22, 8'sd18, 8'sd15, -8'sd4, 8'sd17, 8'sd26, 8'sd22, 8'sd21, 8'sd10, 8'sd10, 8'sd14, 8'sd16, 8'sd25, 8'sd39, 8'sd36, 8'sd42, 8'sd51, 8'sd50, 8'sd40, 8'sd47, 8'sd40, 8'sd21, 8'sd7, 8'sd11, 8'sd14, 8'sd14, 8'sd23, 8'sd20, 8'sd24, 8'sd23, 8'sd36, 8'sd30, 8'sd36, 8'sd38, 8'sd33, 8'sd13, 8'sd11, 8'sd14, 8'sd13, 8'sd12, 8'sd6, 8'sd8, 8'sd21, 8'sd22, 8'sd29, 8'sd31, 8'sd28, 8'sd20, 8'sd7, 8'sd10, 8'sd12, 8'sd11, 8'sd10, 8'sd10, 8'sd12, 8'sd12, 8'sd7, 8'sd10, 8'sd11, 8'sd8, 8'sd12, 8'sd9, 8'sd12, 8'sd14, 8'sd13, 8'sd10,
    8'sd11, 8'sd14, 8'sd14, 8'sd14, 8'sd11, 8'sd12, 8'sd10, 8'sd11, 8'sd14, 8'sd10, 8'sd12, 8'sd13, 8'sd11, 8'sd13, 8'sd12, 8'sd13, 8'sd10, 8'sd12, 8'sd9, 8'sd10, 8'sd18, 8'sd14, 8'sd6, 8'sd3, 8'sd7, 8'sd4, 8'sd10, 8'sd13, 8'sd12, 8'sd13, 8'sd12, 8'sd16, 8'sd20, 8'sd26, 8'sd25, 8'sd26, 8'sd36, 8'sd31, 8'sd10, 8'sd1, 8'sd14, 8'sd14, 8'sd14, 8'sd12, 8'sd20, 8'sd24, 8'sd15, 8'sd17, 8'sd21, 8'sd12, 8'sd11, 8'sd31, 8'sd27, 8'sd24, 8'sd22, 8'sd13, 8'sd13, 8'sd10, 8'sd18, 8'sd18, 8'sd18, 8'sd34, 8'sd32, 8'sd19, 8'sd18, 8'sd26, 8'sd25, 8'sd34, 8'sd35, 8'sd18, 8'sd13, 8'sd12, 8'sd14, 8'sd11, 8'sd4, 8'sd7, 8'sd17, 8'sd17, 8'sd0, 8'sd14, 8'sd14, 8'sd19, 8'sd32, 8'sd12, 8'sd12, 8'sd14, 8'sd6, 8'sd5, 8'sd4, -8'sd2, 8'sd30, 8'sd16, 8'sd3, 8'sd13, -8'sd4, -8'sd12, 8'sd2, 8'sd13, 8'sd10, 8'sd12, 8'sd11, 8'sd7, 8'sd14, 8'sd3, 8'sd21, 8'sd8, -8'sd4, -8'sd3, -8'sd6, 8'sd2, 8'sd9, 8'sd16, 8'sd12, 8'sd16, 8'sd21, -8'sd2, 8'sd4, 8'sd10, 8'sd14, 8'sd0, 8'sd5, 8'sd10, 8'sd19, 8'sd27, 8'sd20, 8'sd12, 8'sd12, 8'sd15, 8'sd30, 8'sd17, 8'sd16, 8'sd17, 8'sd0, 8'sd25, 8'sd27, 8'sd26, 8'sd26, 8'sd39, 8'sd23, 8'sd14, 8'sd11, 8'sd15, 8'sd27, 8'sd37, 8'sd19, 8'sd16, 8'sd5, 8'sd16, 8'sd19, 8'sd17, 8'sd33, 8'sd33, 8'sd16, 8'sd12, 8'sd10, 8'sd16, 8'sd20, 8'sd29, 8'sd13, 8'sd16, 8'sd14, 8'sd7, 8'sd21, 8'sd17, 8'sd15, 8'sd17, 8'sd15, 8'sd13, 8'sd10, 8'sd14, 8'sd9, 8'sd5, 8'sd18, 8'sd20, 8'sd24, 8'sd21, 8'sd22, 8'sd14, 8'sd5, 8'sd12, 8'sd12, 8'sd14, 8'sd13, 8'sd12, 8'sd11, 8'sd12, 8'sd12, 8'sd13, 8'sd16, 8'sd18, 8'sd19, 8'sd11, 8'sd9, 8'sd12, 8'sd12, 8'sd13,
    8'sd17, 8'sd13, 8'sd15, 8'sd17, 8'sd13, 8'sd14, 8'sd17, 8'sd16, 8'sd15, 8'sd13, 8'sd14, 8'sd12, 8'sd12, 8'sd12, 8'sd17, 8'sd16, 8'sd16, 8'sd15, 8'sd19, 8'sd21, 8'sd26, 8'sd21, 8'sd23, 8'sd19, 8'sd14, 8'sd12, 8'sd16, 8'sd14, 8'sd16, 8'sd17, 8'sd20, 8'sd29, 8'sd36, 8'sd26, 8'sd19, 8'sd19, 8'sd20, 8'sd21, 8'sd10, 8'sd10, 8'sd13, 8'sd16, 8'sd16, 8'sd15, 8'sd28, 8'sd36, 8'sd23, 8'sd15, 8'sd23, 8'sd11, 8'sd14, 8'sd15, 8'sd9, 8'sd4, 8'sd2, 8'sd13, 8'sd16, 8'sd18, 8'sd32, 8'sd8, 8'sd0, 8'sd0, 8'sd8, 8'sd23, 8'sd33, 8'sd14, 8'sd13, 8'sd4, -8'sd9, 8'sd9, 8'sd12, 8'sd18, 8'sd6, -8'sd30, -8'sd19, -8'sd15, -8'sd5, -8'sd10, 8'sd27, 8'sd19, 8'sd22, 8'sd16, 8'sd3, 8'sd11, 8'sd16, 8'sd14, -8'sd1, 8'sd4, 8'sd15, 8'sd12, 8'sd15, -8'sd10, 8'sd18, -8'sd2, 8'sd0, 8'sd36, 8'sd34, 8'sd14, 8'sd14, 8'sd15, 8'sd25, 8'sd32, 8'sd25, 8'sd17, 8'sd7, -8'sd11, 8'sd16, 8'sd10, 8'sd24, 8'sd35, 8'sd26, 8'sd15, 8'sd12, 8'sd17, 8'sd17, 8'sd28, 8'sd29, 8'sd16, 8'sd9, 8'sd8, 8'sd30, 8'sd31, 8'sd30, 8'sd32, 8'sd12, 8'sd12, 8'sd14, 8'sd22, 8'sd13, 8'sd16, 8'sd16, 8'sd18, 8'sd8, 8'sd23, 8'sd30, 8'sd26, 8'sd25, 8'sd18, 8'sd12, 8'sd17, 8'sd16, 8'sd21, 8'sd19, 8'sd23, 8'sd17, 8'sd22, 8'sd23, 8'sd18, 8'sd20, 8'sd22, 8'sd21, 8'sd3, 8'sd13, 8'sd15, 8'sd13, 8'sd19, 8'sd16, 8'sd18, 8'sd16, 8'sd21, 8'sd15, 8'sd17, 8'sd7, 8'sd10, 8'sd5, 8'sd9, 8'sd13, 8'sd12, 8'sd14, 8'sd16, 8'sd22, 8'sd25, 8'sd25, 8'sd22, 8'sd19, 8'sd14, 8'sd15, 8'sd0, 8'sd2, 8'sd11, 8'sd16, 8'sd17, 8'sd12, 8'sd17, 8'sd13, 8'sd14, 8'sd17, 8'sd15, 8'sd15, 8'sd16, 8'sd13, 8'sd16, 8'sd15, 8'sd14, 8'sd15, 8'sd14,
    8'sd15, 8'sd15, 8'sd16, 8'sd15, 8'sd15, 8'sd17, 8'sd15, 8'sd15, 8'sd17, 8'sd15, 8'sd19, 8'sd16, 8'sd15, 8'sd16, 8'sd15, 8'sd18, 8'sd19, 8'sd15, 8'sd15, 8'sd16, 8'sd13, 8'sd14, 8'sd15, 8'sd17, 8'sd18, 8'sd15, 8'sd18, 8'sd16, 8'sd17, 8'sd15, 8'sd20, 8'sd17, 8'sd13, 8'sd22, 8'sd16, 8'sd13, 8'sd15, 8'sd13, 8'sd16, 8'sd24, 8'sd22, 8'sd18, 8'sd18, 8'sd18, 8'sd23, 8'sd13, 8'sd20, 8'sd18, 8'sd20, 8'sd18, 8'sd21, 8'sd18, 8'sd20, 8'sd18, 8'sd30, 8'sd21, 8'sd18, 8'sd21, 8'sd20, 8'sd16, 8'sd25, 8'sd19, 8'sd19, 8'sd14, 8'sd13, 8'sd10, 8'sd11, 8'sd13, 8'sd29, 8'sd20, 8'sd19, 8'sd22, 8'sd13, 8'sd7, 8'sd6, 8'sd4, 8'sd13, -8'sd1, 8'sd2, 8'sd6, 8'sd0, -8'sd5, 8'sd11, 8'sd17, 8'sd19, 8'sd22, 8'sd17, 8'sd9, 8'sd16, 8'sd15, 8'sd22, 8'sd14, 8'sd16, 8'sd12, 8'sd4, -8'sd4, 8'sd3, 8'sd15, 8'sd16, 8'sd16, 8'sd13, 8'sd6, 8'sd24, 8'sd22, 8'sd23, 8'sd17, 8'sd5, 8'sd9, 8'sd16, 8'sd24, 8'sd14, 8'sd16, 8'sd19, 8'sd20, -8'sd6, -8'sd37, -8'sd24, 8'sd10, 8'sd28, 8'sd4, 8'sd10, 8'sd24, 8'sd18, 8'sd26, 8'sd20, 8'sd17, 8'sd18, 8'sd25, 8'sd1, -8'sd18, -8'sd36, -8'sd62, -8'sd55, -8'sd5, 8'sd14, 8'sd17, 8'sd17, 8'sd19, 8'sd17, 8'sd17, 8'sd18, 8'sd23, 8'sd22, 8'sd14, 8'sd23, 8'sd33, 8'sd32, 8'sd20, 8'sd8, 8'sd11, 8'sd16, 8'sd12, 8'sd16, 8'sd15, 8'sd16, 8'sd18, 8'sd28, 8'sd27, 8'sd23, 8'sd30, 8'sd28, 8'sd28, 8'sd19, 8'sd18, 8'sd9, 8'sd15, 8'sd15, 8'sd18, 8'sd16, 8'sd17, 8'sd24, 8'sd41, 8'sd37, 8'sd30, 8'sd24, 8'sd19, 8'sd17, 8'sd11, 8'sd16, 8'sd21, 8'sd14, 8'sd14, 8'sd16, 8'sd15, 8'sd16, 8'sd17, 8'sd16, 8'sd20, 8'sd17, 8'sd22, 8'sd20, 8'sd18, 8'sd16, 8'sd17, 8'sd15, 8'sd19,
    8'sd10, 8'sd12, 8'sd11, 8'sd11, 8'sd11, 8'sd12, 8'sd12, 8'sd13, 8'sd14, 8'sd11, 8'sd11, 8'sd12, 8'sd15, 8'sd12, 8'sd10, 8'sd14, 8'sd13, 8'sd12, 8'sd11, 8'sd11, 8'sd11, 8'sd13, 8'sd13, 8'sd17, 8'sd17, 8'sd13, 8'sd14, 8'sd12, 8'sd11, 8'sd11, 8'sd15, 8'sd14, 8'sd17, 8'sd15, 8'sd9, 8'sd4, 8'sd8, 8'sd19, 8'sd17, 8'sd17, 8'sd16, 8'sd13, 8'sd12, 8'sd11, 8'sd19, 8'sd19, 8'sd21, 8'sd19, 8'sd16, 8'sd13, 8'sd15, 8'sd29, 8'sd15, 8'sd14, 8'sd18, 8'sd12, 8'sd12, 8'sd14, 8'sd16, 8'sd18, 8'sd11, 8'sd14, 8'sd9, 8'sd11, 8'sd12, 8'sd14, 8'sd28, 8'sd25, 8'sd25, 8'sd15, 8'sd10, 8'sd12, 8'sd16, 8'sd17, 8'sd9, 8'sd13, 8'sd14, 8'sd13, 8'sd32, 8'sd4, -8'sd3, 8'sd2, 8'sd8, 8'sd14, 8'sd12, 8'sd15, 8'sd27, 8'sd23, 8'sd19, 8'sd22, 8'sd13, 8'sd20, 8'sd37, 8'sd28, 8'sd10, -8'sd8, -8'sd2, 8'sd10, 8'sd14, 8'sd14, 8'sd15, 8'sd4, -8'sd7, -8'sd2, 8'sd4, 8'sd27, 8'sd27, 8'sd24, 8'sd29, 8'sd16, 8'sd5, 8'sd11, 8'sd12, 8'sd15, 8'sd5, 8'sd5, 8'sd0, -8'sd26, 8'sd15, 8'sd33, 8'sd14, 8'sd25, 8'sd20, 8'sd6, 8'sd4, 8'sd11, 8'sd12, 8'sd19, 8'sd15, 8'sd15, 8'sd2, -8'sd21, 8'sd33, 8'sd29, 8'sd24, 8'sd23, 8'sd16, -8'sd2, 8'sd1, 8'sd13, 8'sd14, 8'sd12, 8'sd13, 8'sd2, -8'sd3, -8'sd4, 8'sd15, 8'sd26, 8'sd41, 8'sd22, 8'sd15, 8'sd9, 8'sd10, 8'sd11, 8'sd12, 8'sd11, 8'sd15, -8'sd4, -8'sd2, 8'sd6, -8'sd3, 8'sd15, 8'sd23, 8'sd22, 8'sd18, 8'sd17, 8'sd15, 8'sd13, 8'sd11, 8'sd14, 8'sd23, 8'sd34, 8'sd24, 8'sd12, 8'sd10, 8'sd18, 8'sd22, 8'sd23, 8'sd23, 8'sd19, 8'sd10, 8'sd12, 8'sd11, 8'sd14, 8'sd13, 8'sd16, 8'sd18, 8'sd16, 8'sd18, 8'sd17, 8'sd15, 8'sd14, 8'sd14, 8'sd14, 8'sd12, 8'sd13,
    8'sd20, 8'sd19, 8'sd19, 8'sd19, 8'sd16, 8'sd17, 8'sd16, 8'sd20, 8'sd16, 8'sd16, 8'sd19, 8'sd20, 8'sd16, 8'sd20, 8'sd18, 8'sd19, 8'sd17, 8'sd19, 8'sd23, 8'sd26, 8'sd24, 8'sd17, 8'sd16, 8'sd13, 8'sd11, 8'sd16, 8'sd15, 8'sd18, 8'sd18, 8'sd17, 8'sd20, 8'sd19, 8'sd15, 8'sd17, 8'sd15, 8'sd16, 8'sd24, 8'sd12, 8'sd10, 8'sd8, 8'sd16, 8'sd20, 8'sd20, 8'sd18, 8'sd13, 8'sd1, 8'sd6, 8'sd14, 8'sd7, 8'sd20, 8'sd20, 8'sd16, 8'sd17, 8'sd10, 8'sd4, 8'sd18, 8'sd17, 8'sd16, 8'sd13, 8'sd10, 8'sd17, 8'sd25, 8'sd6, 8'sd9, 8'sd16, 8'sd9, 8'sd8, -8'sd3, -8'sd3, 8'sd20, 8'sd17, 8'sd16, 8'sd9, -8'sd2, 8'sd6, -8'sd2, -8'sd12, 8'sd6, 8'sd26, 8'sd6, 8'sd12, -8'sd4, 8'sd13, 8'sd18, 8'sd19, 8'sd18, -8'sd9, -8'sd33, -8'sd27, -8'sd13, 8'sd1, 8'sd1, 8'sd7, 8'sd7, 8'sd16, 8'sd0, 8'sd14, 8'sd21, 8'sd18, 8'sd20, 8'sd5, 8'sd13, 8'sd28, 8'sd30, 8'sd29, 8'sd10, 8'sd5, -8'sd10, -8'sd10, 8'sd4, 8'sd24, 8'sd24, 8'sd17, 8'sd19, 8'sd28, 8'sd29, 8'sd23, 8'sd22, 8'sd42, 8'sd16, -8'sd2, 8'sd0, 8'sd18, 8'sd27, 8'sd38, 8'sd23, 8'sd18, 8'sd15, 8'sd25, 8'sd22, 8'sd29, 8'sd29, 8'sd41, -8'sd15, 8'sd1, 8'sd12, 8'sd22, 8'sd25, 8'sd39, 8'sd22, 8'sd17, 8'sd18, 8'sd27, 8'sd16, 8'sd22, 8'sd24, 8'sd7, 8'sd0, 8'sd10, 8'sd22, 8'sd8, 8'sd23, 8'sd28, 8'sd19, 8'sd18, 8'sd17, 8'sd26, 8'sd14, 8'sd12, 8'sd8, 8'sd15, 8'sd6, 8'sd10, 8'sd26, 8'sd22, 8'sd21, 8'sd19, 8'sd19, 8'sd20, 8'sd17, 8'sd13, 8'sd2, -8'sd2, 8'sd3, 8'sd14, 8'sd13, 8'sd11, 8'sd9, 8'sd16, 8'sd17, 8'sd20, 8'sd21, 8'sd20, 8'sd19, 8'sd21, 8'sd15, 8'sd17, 8'sd17, 8'sd16, 8'sd15, 8'sd16, 8'sd15, 8'sd16, 8'sd20, 8'sd17, 8'sd18,
    8'sd20, 8'sd18, 8'sd19, 8'sd16, 8'sd20, 8'sd16, 8'sd18, 8'sd16, 8'sd16, 8'sd20, 8'sd17, 8'sd18, 8'sd19, 8'sd21, 8'sd20, 8'sd20, 8'sd18, 8'sd16, 8'sd15, 8'sd10, 8'sd7, 8'sd2, 8'sd5, 8'sd13, 8'sd12, 8'sd15, 8'sd18, 8'sd18, 8'sd17, 8'sd21, 8'sd17, 8'sd7, -8'sd2, -8'sd5, -8'sd3, 8'sd0, -8'sd7, -8'sd6, 8'sd1, 8'sd10, 8'sd14, 8'sd19, 8'sd21, 8'sd19, 8'sd21, 8'sd11, 8'sd9, 8'sd8, 8'sd3, 8'sd14, 8'sd17, 8'sd14, 8'sd21, 8'sd26, 8'sd28, 8'sd19, 8'sd18, 8'sd25, 8'sd22, 8'sd17, 8'sd17, -8'sd5, 8'sd21, 8'sd21, 8'sd33, 8'sd28, 8'sd23, 8'sd26, 8'sd32, 8'sd22, 8'sd17, 8'sd23, 8'sd12, 8'sd1, 8'sd14, 8'sd32, 8'sd18, 8'sd20, 8'sd22, 8'sd13, 8'sd17, 8'sd30, 8'sd35, 8'sd22, 8'sd21, 8'sd22, 8'sd18, 8'sd31, 8'sd33, 8'sd25, 8'sd1, 8'sd18, 8'sd16, 8'sd2, -8'sd2, -8'sd4, 8'sd11, 8'sd19, 8'sd18, 8'sd22, 8'sd16, 8'sd17, 8'sd22, 8'sd6, 8'sd8, 8'sd16, 8'sd37, 8'sd14, 8'sd14, 8'sd7, 8'sd10, 8'sd19, 8'sd17, 8'sd13, -8'sd1, 8'sd5, 8'sd20, 8'sd18, 8'sd23, 8'sd21, 8'sd11, 8'sd6, 8'sd12, -8'sd4, 8'sd1, 8'sd15, 8'sd19, 8'sd14, -8'sd14, -8'sd5, 8'sd6, 8'sd13, 8'sd27, 8'sd14, -8'sd5, 8'sd5, 8'sd1, -8'sd16, 8'sd2, 8'sd19, 8'sd18, 8'sd14, -8'sd12, -8'sd4, 8'sd2, -8'sd4, 8'sd4, 8'sd11, 8'sd2, -8'sd2, -8'sd1, 8'sd5, 8'sd12, 8'sd17, 8'sd17, 8'sd15, 8'sd13, 8'sd14, 8'sd15, 8'sd16, 8'sd10, 8'sd12, 8'sd8, 8'sd4, 8'sd1, 8'sd17, 8'sd18, 8'sd20, 8'sd20, 8'sd21, 8'sd17, 8'sd21, 8'sd17, 8'sd13, 8'sd10, 8'sd17, 8'sd10, 8'sd18, 8'sd17, 8'sd21, 8'sd16, 8'sd20, 8'sd17, 8'sd17, 8'sd21, 8'sd20, 8'sd19, 8'sd20, 8'sd20, 8'sd23, 8'sd17, 8'sd19, 8'sd17, 8'sd20, 8'sd17, 8'sd18,
    8'sd15, 8'sd17, 8'sd17, 8'sd19, 8'sd17, 8'sd20, 8'sd20, 8'sd19, 8'sd17, 8'sd16, 8'sd16, 8'sd17, 8'sd16, 8'sd19, 8'sd17, 8'sd17, 8'sd18, 8'sd17, 8'sd24, 8'sd22, 8'sd21, 8'sd26, 8'sd19, 8'sd17, 8'sd13, 8'sd16, 8'sd17, 8'sd19, 8'sd19, 8'sd19, 8'sd16, 8'sd18, 8'sd15, 8'sd14, 8'sd24, 8'sd24, 8'sd5, 8'sd3, 8'sd10, 8'sd13, 8'sd15, 8'sd17, 8'sd18, 8'sd19, 8'sd16, 8'sd25, 8'sd13, 8'sd14, 8'sd5, -8'sd12, 8'sd9, 8'sd10, 8'sd7, 8'sd4, 8'sd10, 8'sd14, 8'sd20, 8'sd26, 8'sd25, 8'sd23, 8'sd15, 8'sd18, 8'sd11, 8'sd10, 8'sd8, 8'sd12, 8'sd11, 8'sd14, 8'sd7, 8'sd15, 8'sd18, 8'sd28, 8'sd27, 8'sd18, 8'sd18, 8'sd27, 8'sd13, 8'sd8, 8'sd13, 8'sd13, 8'sd18, 8'sd16, 8'sd13, 8'sd14, 8'sd18, 8'sd27, 8'sd26, 8'sd25, 8'sd29, 8'sd11, -8'sd29, 8'sd10, 8'sd6, 8'sd16, 8'sd12, 8'sd19, 8'sd21, 8'sd16, 8'sd16, 8'sd19, 8'sd11, 8'sd14, 8'sd5, -8'sd33, 8'sd1, 8'sd21, 8'sd6, 8'sd13, 8'sd14, 8'sd29, 8'sd22, 8'sd16, 8'sd15, 8'sd14, 8'sd6, 8'sd2, -8'sd27, -8'sd35, 8'sd34, 8'sd30, 8'sd21, 8'sd14, 8'sd18, 8'sd14, 8'sd24, 8'sd16, 8'sd19, 8'sd16, 8'sd4, -8'sd11, -8'sd22, -8'sd3, 8'sd59, 8'sd30, 8'sd20, 8'sd20, 8'sd6, 8'sd8, 8'sd17, 8'sd16, 8'sd19, 8'sd16, 8'sd2, -8'sd3, -8'sd4, 8'sd22, 8'sd36, 8'sd36, 8'sd23, 8'sd21, 8'sd2, 8'sd10, 8'sd18, 8'sd20, 8'sd16, 8'sd17, 8'sd13, 8'sd10, 8'sd6, -8'sd4, 8'sd8, 8'sd16, 8'sd27, 8'sd25, 8'sd8, 8'sd9, 8'sd18, 8'sd18, 8'sd16, 8'sd16, 8'sd15, 8'sd11, 8'sd10, 8'sd5, 8'sd15, 8'sd15, 8'sd14, 8'sd14, 8'sd12, 8'sd13, 8'sd17, 8'sd15, 8'sd19, 8'sd16, 8'sd17, 8'sd15, 8'sd20, 8'sd16, 8'sd14, 8'sd16, 8'sd18, 8'sd25, 8'sd20, 8'sd19, 8'sd17, 8'sd17,
    8'sd15, 8'sd13, 8'sd13, 8'sd11, 8'sd11, 8'sd12, 8'sd14, 8'sd14, 8'sd14, 8'sd14, 8'sd13, 8'sd11, 8'sd16, 8'sd12, 8'sd14, 8'sd15, 8'sd14, 8'sd7, -8'sd1, 8'sd2, -8'sd2, 8'sd9, 8'sd20, 8'sd15, 8'sd11, 8'sd11, 8'sd12, 8'sd14, 8'sd16, 8'sd16, 8'sd17, 8'sd11, 8'sd12, 8'sd13, 8'sd19, 8'sd3, -8'sd1, 8'sd1, 8'sd18, 8'sd25, 8'sd21, 8'sd17, 8'sd12, 8'sd13, 8'sd22, 8'sd20, 8'sd24, 8'sd25, 8'sd23, 8'sd27, 8'sd29, 8'sd28, 8'sd29, 8'sd41, 8'sd21, 8'sd13, 8'sd15, 8'sd18, 8'sd16, 8'sd17, 8'sd20, 8'sd16, 8'sd29, 8'sd31, 8'sd48, 8'sd37, 8'sd26, 8'sd28, 8'sd13, 8'sd10, 8'sd15, 8'sd17, 8'sd14, 8'sd19, 8'sd23, 8'sd25, 8'sd21, 8'sd8, 8'sd15, 8'sd12, 8'sd24, 8'sd18, 8'sd13, 8'sd17, 8'sd15, 8'sd15, 8'sd25, 8'sd43, 8'sd39, 8'sd34, 8'sd20, 8'sd3, 8'sd11, 8'sd18, 8'sd14, 8'sd22, 8'sd14, 8'sd15, 8'sd15, 8'sd12, 8'sd30, 8'sd22, 8'sd24, 8'sd20, 8'sd5, 8'sd7, 8'sd16, 8'sd18, 8'sd8, 8'sd14, 8'sd8, 8'sd12, 8'sd12, 8'sd10, 8'sd3, 8'sd8, 8'sd23, 8'sd16, 8'sd18, 8'sd5, 8'sd22, 8'sd17, 8'sd14, 8'sd18, 8'sd2, 8'sd13, 8'sd16, 8'sd11, -8'sd2, 8'sd6, -8'sd1, 8'sd0, -8'sd1, -8'sd3, 8'sd10, 8'sd13, 8'sd8, 8'sd8, -8'sd2, 8'sd15, 8'sd15, 8'sd13, 8'sd0, -8'sd3, -8'sd8, -8'sd9, -8'sd3, -8'sd1, 8'sd7, 8'sd2, 8'sd16, 8'sd0, 8'sd4, 8'sd11, 8'sd14, 8'sd14, 8'sd9, 8'sd21, 8'sd15, 8'sd19, 8'sd26, 8'sd20, 8'sd17, 8'sd10, 8'sd17, 8'sd9, 8'sd11, 8'sd15, 8'sd14, 8'sd15, 8'sd19, 8'sd27, 8'sd30, 8'sd37, 8'sd36, 8'sd37, 8'sd29, 8'sd17, 8'sd16, 8'sd15, 8'sd15, 8'sd14, 8'sd13, 8'sd12, 8'sd12, 8'sd16, 8'sd13, 8'sd16, 8'sd18, 8'sd19, 8'sd13, 8'sd15, 8'sd15, 8'sd16, 8'sd14, 8'sd15,
    8'sd16, 8'sd18, 8'sd16, 8'sd14, 8'sd16, 8'sd14, 8'sd16, 8'sd18, 8'sd15, 8'sd14, 8'sd16, 8'sd16, 8'sd15, 8'sd18, 8'sd17, 8'sd15, 8'sd16, 8'sd16, 8'sd15, 8'sd22, 8'sd31, 8'sd28, 8'sd18, 8'sd4, 8'sd5, 8'sd7, 8'sd16, 8'sd15, 8'sd16, 8'sd14, 8'sd17, 8'sd24, 8'sd25, 8'sd32, 8'sd36, 8'sd30, 8'sd14, 8'sd12, 8'sd0, 8'sd1, 8'sd18, 8'sd15, 8'sd15, 8'sd15, 8'sd19, 8'sd9, 8'sd5, 8'sd19, 8'sd36, 8'sd31, 8'sd27, 8'sd12, 8'sd28, 8'sd22, 8'sd22, 8'sd19, 8'sd18, 8'sd15, 8'sd16, 8'sd12, 8'sd7, 8'sd0, 8'sd27, 8'sd41, 8'sd23, 8'sd17, 8'sd26, 8'sd29, 8'sd22, 8'sd14, 8'sd14, 8'sd16, 8'sd15, -8'sd1, -8'sd7, -8'sd27, -8'sd17, 8'sd31, 8'sd24, 8'sd20, 8'sd5, 8'sd3, 8'sd20, 8'sd14, 8'sd13, 8'sd14, -8'sd7, -8'sd30, -8'sd6, -8'sd3, -8'sd7, 8'sd24, 8'sd5, 8'sd11, 8'sd5, -8'sd7, 8'sd15, 8'sd18, 8'sd17, 8'sd15, 8'sd10, 8'sd10, 8'sd16, 8'sd10, 8'sd17, 8'sd27, 8'sd10, 8'sd12, 8'sd4, 8'sd2, 8'sd21, 8'sd20, 8'sd17, 8'sd22, 8'sd34, 8'sd10, 8'sd4, -8'sd4, 8'sd1, 8'sd16, 8'sd5, 8'sd9, 8'sd7, 8'sd7, 8'sd24, 8'sd17, 8'sd17, 8'sd20, 8'sd41, 8'sd25, 8'sd23, 8'sd5, 8'sd14, 8'sd23, 8'sd18, 8'sd25, 8'sd17, 8'sd23, 8'sd32, 8'sd15, 8'sd16, 8'sd20, 8'sd33, 8'sd37, 8'sd29, 8'sd25, 8'sd16, 8'sd17, 8'sd20, 8'sd22, 8'sd24, 8'sd25, 8'sd22, 8'sd14, 8'sd14, 8'sd16, 8'sd17, 8'sd22, 8'sd24, 8'sd23, 8'sd4, 8'sd8, 8'sd12, 8'sd20, 8'sd17, 8'sd21, 8'sd20, 8'sd18, 8'sd15, 8'sd19, 8'sd17, 8'sd12, 8'sd12, 8'sd13, 8'sd22, 8'sd12, 8'sd8, 8'sd4, 8'sd6, 8'sd14, 8'sd19, 8'sd16, 8'sd14, 8'sd15, 8'sd14, 8'sd16, 8'sd13, 8'sd13, 8'sd14, 8'sd14, 8'sd13, 8'sd17, 8'sd14, 8'sd14, 8'sd17, 8'sd14,
    8'sd16, 8'sd15, 8'sd13, 8'sd13, 8'sd13, 8'sd14, 8'sd14, 8'sd13, 8'sd12, 8'sd12, 8'sd12, 8'sd14, 8'sd14, 8'sd13, 8'sd14, 8'sd14, 8'sd16, 8'sd11, 8'sd11, 8'sd10, 8'sd11, 8'sd14, 8'sd24, 8'sd23, 8'sd18, 8'sd13, 8'sd16, 8'sd13, 8'sd14, 8'sd16, 8'sd15, 8'sd9, 8'sd13, 8'sd9, 8'sd13, 8'sd20, 8'sd37, 8'sd35, 8'sd32, 8'sd27, 8'sd16, 8'sd15, 8'sd16, 8'sd11, 8'sd12, 8'sd17, 8'sd25, -8'sd7, -8'sd15, -8'sd9, -8'sd4, 8'sd3, 8'sd6, 8'sd41, 8'sd24, 8'sd15, 8'sd16, 8'sd11, 8'sd7, 8'sd4, 8'sd6, -8'sd5, -8'sd21, -8'sd19, 8'sd4, -8'sd1, 8'sd10, 8'sd17, 8'sd33, 8'sd15, 8'sd16, 8'sd11, -8'sd1, -8'sd6, 8'sd8, 8'sd14, -8'sd1, 8'sd15, 8'sd17, 8'sd0, 8'sd1, 8'sd7, 8'sd20, 8'sd14, 8'sd15, 8'sd13, 8'sd11, 8'sd26, 8'sd20, 8'sd57, 8'sd28, -8'sd2, -8'sd4, 8'sd2, 8'sd7, 8'sd25, 8'sd15, 8'sd12, 8'sd16, 8'sd14, 8'sd30, 8'sd33, 8'sd48, 8'sd43, 8'sd15, 8'sd6, 8'sd24, 8'sd21, 8'sd20, 8'sd38, 8'sd22, 8'sd12, 8'sd16, 8'sd18, 8'sd24, 8'sd35, 8'sd20, 8'sd6, 8'sd14, 8'sd26, 8'sd28, 8'sd26, 8'sd30, 8'sd31, 8'sd17, 8'sd12, 8'sd16, 8'sd14, 8'sd31, 8'sd34, 8'sd3, 8'sd1, 8'sd18, 8'sd29, 8'sd24, 8'sd14, 8'sd18, 8'sd20, 8'sd11, 8'sd11, 8'sd16, 8'sd16, 8'sd23, 8'sd22, 8'sd23, 8'sd26, 8'sd29, 8'sd29, 8'sd23, 8'sd19, 8'sd13, 8'sd15, 8'sd12, 8'sd16, 8'sd13, 8'sd12, 8'sd12, 8'sd11, 8'sd9, 8'sd13, 8'sd13, 8'sd8, 8'sd14, 8'sd22, 8'sd14, 8'sd3, 8'sd14, 8'sd13, 8'sd15, 8'sd13, 8'sd12, -8'sd1, -8'sd14, -8'sd6, -8'sd2, 8'sd8, 8'sd8, 8'sd6, 8'sd4, 8'sd9, 8'sd13, 8'sd15, 8'sd15, 8'sd12, 8'sd14, 8'sd7, 8'sd7, 8'sd2, -8'sd1, -8'sd6, -8'sd1, 8'sd1, 8'sd12, 8'sd12, 8'sd14, 8'sd12,
    8'sd15, 8'sd12, 8'sd15, 8'sd16, 8'sd12, 8'sd14, 8'sd13, 8'sd17, 8'sd14, 8'sd16, 8'sd13, 8'sd15, 8'sd17, 8'sd15, 8'sd14, 8'sd14, 8'sd16, 8'sd16, 8'sd15, 8'sd14, 8'sd10, 8'sd8, 8'sd9, 8'sd10, 8'sd7, 8'sd12, 8'sd16, 8'sd16, 8'sd16, 8'sd16, 8'sd13, 8'sd13, 8'sd13, 8'sd15, 8'sd18, 8'sd14, 8'sd18, 8'sd20, 8'sd14, 8'sd6, 8'sd16, 8'sd15, 8'sd14, 8'sd15, 8'sd15, 8'sd14, 8'sd22, 8'sd24, 8'sd17, 8'sd3, 8'sd26, 8'sd34, 8'sd17, 8'sd5, 8'sd12, 8'sd17, 8'sd15, 8'sd12, 8'sd20, 8'sd31, 8'sd25, 8'sd24, 8'sd14, 8'sd8, 8'sd36, 8'sd28, 8'sd18, 8'sd13, 8'sd4, 8'sd16, 8'sd17, 8'sd15, 8'sd25, 8'sd27, 8'sd15, 8'sd13, -8'sd22, 8'sd27, 8'sd36, 8'sd11, 8'sd12, 8'sd15, 8'sd9, 8'sd16, 8'sd14, 8'sd13, 8'sd18, -8'sd5, -8'sd13, -8'sd26, -8'sd2, 8'sd50, 8'sd19, 8'sd28, 8'sd43, 8'sd15, 8'sd17, 8'sd16, 8'sd13, 8'sd13, 8'sd4, -8'sd13, -8'sd7, 8'sd16, 8'sd39, 8'sd36, 8'sd28, 8'sd31, 8'sd11, -8'sd10, 8'sd10, 8'sd14, 8'sd17, 8'sd11, 8'sd5, 8'sd11, 8'sd28, 8'sd23, 8'sd36, 8'sd32, 8'sd25, 8'sd6, 8'sd0, -8'sd5, 8'sd14, 8'sd13, 8'sd15, 8'sd12, -8'sd3, 8'sd0, 8'sd8, 8'sd0, 8'sd17, 8'sd12, 8'sd0, 8'sd6, 8'sd9, 8'sd10, 8'sd18, 8'sd13, 8'sd13, 8'sd15, 8'sd19, 8'sd15, 8'sd11, 8'sd1, 8'sd1, 8'sd8, 8'sd6, 8'sd5, 8'sd18, 8'sd18, 8'sd17, 8'sd12, 8'sd17, 8'sd16, 8'sd23, 8'sd24, 8'sd14, 8'sd8, 8'sd11, 8'sd13, 8'sd7, 8'sd9, 8'sd22, 8'sd21, 8'sd18, 8'sd12, 8'sd14, 8'sd15, 8'sd17, 8'sd20, 8'sd14, 8'sd6, 8'sd12, 8'sd14, 8'sd12, 8'sd17, 8'sd23, 8'sd18, 8'sd17, 8'sd14, 8'sd14, 8'sd15, 8'sd18, 8'sd15, 8'sd19, 8'sd18, 8'sd20, 8'sd23, 8'sd15, 8'sd14, 8'sd15, 8'sd16, 8'sd17, 8'sd12,
    8'sd16, 8'sd13, 8'sd14, 8'sd13, 8'sd15, 8'sd12, 8'sd13, 8'sd13, 8'sd16, 8'sd15, 8'sd12, 8'sd15, 8'sd16, 8'sd11, 8'sd16, 8'sd16, 8'sd15, 8'sd16, 8'sd23, 8'sd28, 8'sd34, 8'sd34, 8'sd26, 8'sd24, 8'sd19, 8'sd20, 8'sd15, 8'sd16, 8'sd14, 8'sd15, 8'sd17, 8'sd19, 8'sd17, 8'sd10, 8'sd20, 8'sd23, 8'sd10, 8'sd5, 8'sd19, 8'sd15, 8'sd16, 8'sd12, 8'sd15, 8'sd14, 8'sd15, 8'sd0, 8'sd7, 8'sd0, 8'sd9, 8'sd40, 8'sd30, -8'sd8, 8'sd4, -8'sd8, 8'sd7, 8'sd13, 8'sd11, 8'sd12, 8'sd15, 8'sd17, 8'sd13, -8'sd1, 8'sd2, 8'sd49, 8'sd3, -8'sd5, 8'sd15, -8'sd14, -8'sd12, 8'sd14, 8'sd12, 8'sd17, 8'sd18, 8'sd18, -8'sd2, -8'sd8, -8'sd17, 8'sd65, 8'sd7, 8'sd11, 8'sd9, 8'sd10, 8'sd6, 8'sd14, 8'sd12, 8'sd16, 8'sd20, 8'sd5, 8'sd19, 8'sd6, -8'sd14, 8'sd56, 8'sd20, 8'sd21, 8'sd10, 8'sd30, 8'sd21, 8'sd15, 8'sd12, 8'sd18, 8'sd5, 8'sd17, 8'sd12, 8'sd7, 8'sd15, 8'sd39, 8'sd21, 8'sd16, 8'sd22, 8'sd13, 8'sd18, 8'sd12, 8'sd15, 8'sd19, 8'sd11, 8'sd26, 8'sd17, 8'sd16, 8'sd22, 8'sd30, 8'sd17, 8'sd16, 8'sd14, 8'sd6, 8'sd12, 8'sd13, 8'sd13, 8'sd18, 8'sd10, 8'sd4, 8'sd11, 8'sd12, 8'sd20, 8'sd23, 8'sd22, 8'sd21, 8'sd14, 8'sd10, 8'sd10, 8'sd13, 8'sd12, 8'sd18, 8'sd18, 8'sd19, 8'sd5, 8'sd3, 8'sd23, 8'sd31, 8'sd22, 8'sd16, 8'sd1, -8'sd2, 8'sd12, 8'sd14, 8'sd13, 8'sd16, 8'sd17, 8'sd6, -8'sd1, -8'sd1, 8'sd2, 8'sd18, 8'sd15, 8'sd9, 8'sd10, 8'sd12, 8'sd15, 8'sd15, 8'sd15, 8'sd14, 8'sd16, 8'sd23, 8'sd20, 8'sd25, 8'sd9, 8'sd12, 8'sd20, 8'sd29, 8'sd33, 8'sd18, 8'sd13, 8'sd14, 8'sd13, 8'sd15, 8'sd15, 8'sd17, 8'sd24, 8'sd24, 8'sd23, 8'sd24, 8'sd20, 8'sd16, 8'sd16, 8'sd16, 8'sd13, 8'sd15,
    8'sd19, 8'sd17, 8'sd19, 8'sd19, 8'sd17, 8'sd18, 8'sd20, 8'sd21, 8'sd19, 8'sd18, 8'sd17, 8'sd17, 8'sd19, 8'sd18, 8'sd16, 8'sd18, 8'sd16, 8'sd20, 8'sd19, 8'sd22, 8'sd24, 8'sd25, 8'sd20, 8'sd23, 8'sd22, 8'sd21, 8'sd18, 8'sd20, 8'sd20, 8'sd18, 8'sd17, 8'sd14, 8'sd4, -8'sd1, 8'sd1, 8'sd2, 8'sd5, 8'sd27, 8'sd22, 8'sd29, 8'sd17, 8'sd16, 8'sd18, 8'sd14, 8'sd11, -8'sd6, -8'sd15, 8'sd6, 8'sd11, 8'sd17, 8'sd5, 8'sd17, 8'sd4, 8'sd8, 8'sd14, 8'sd16, 8'sd19, 8'sd15, -8'sd6, -8'sd20, 8'sd5, 8'sd14, 8'sd14, 8'sd9, 8'sd10, -8'sd5, -8'sd12, 8'sd0, 8'sd10, 8'sd17, 8'sd16, 8'sd11, -8'sd7, 8'sd12, 8'sd29, 8'sd31, 8'sd26, 8'sd14, -8'sd10, 8'sd0, 8'sd8, 8'sd20, 8'sd8, 8'sd16, 8'sd16, 8'sd12, 8'sd17, 8'sd40, 8'sd30, 8'sd14, 8'sd19, 8'sd26, 8'sd18, 8'sd20, 8'sd21, 8'sd44, 8'sd26, 8'sd15, 8'sd16, 8'sd15, 8'sd14, 8'sd35, 8'sd25, 8'sd12, 8'sd8, 8'sd30, 8'sd24, -8'sd1, 8'sd14, 8'sd19, 8'sd14, 8'sd13, 8'sd20, 8'sd13, -8'sd5, 8'sd10, 8'sd28, 8'sd34, 8'sd19, 8'sd31, 8'sd2, 8'sd5, 8'sd1, 8'sd6, 8'sd8, 8'sd17, 8'sd19, 8'sd13, -8'sd3, -8'sd8, -8'sd2, 8'sd13, 8'sd24, 8'sd15, 8'sd5, 8'sd5, 8'sd15, 8'sd12, 8'sd4, 8'sd18, 8'sd15, 8'sd17, 8'sd4, 8'sd8, 8'sd14, 8'sd24, 8'sd25, 8'sd26, 8'sd20, 8'sd10, 8'sd13, 8'sd9, 8'sd15, 8'sd18, 8'sd18, 8'sd16, 8'sd14, 8'sd4, 8'sd26, 8'sd15, 8'sd17, 8'sd13, 8'sd23, 8'sd6, 8'sd7, 8'sd13, 8'sd17, 8'sd16, 8'sd18, 8'sd20, 8'sd21, 8'sd16, 8'sd17, 8'sd10, 8'sd4, 8'sd5, 8'sd13, 8'sd14, 8'sd21, 8'sd22, 8'sd18, 8'sd17, 8'sd19, 8'sd20, 8'sd17, 8'sd21, 8'sd19, 8'sd20, 8'sd21, 8'sd21, 8'sd17, 8'sd15, 8'sd17, 8'sd19, 8'sd17, 8'sd20,
    8'sd10, 8'sd13, 8'sd11, 8'sd9, 8'sd11, 8'sd10, 8'sd11, 8'sd11, 8'sd8, 8'sd11, 8'sd12, 8'sd10, 8'sd11, 8'sd12, 8'sd9, 8'sd13, 8'sd8, 8'sd10, 8'sd12, 8'sd10, -8'sd1, 8'sd0, 8'sd11, 8'sd17, 8'sd14, 8'sd11, 8'sd9, 8'sd11, 8'sd9, 8'sd9, 8'sd8, 8'sd5, 8'sd10, 8'sd8, 8'sd12, 8'sd11, 8'sd21, 8'sd27, 8'sd25, 8'sd22, 8'sd14, 8'sd11, 8'sd10, 8'sd10, 8'sd4, 8'sd16, 8'sd16, 8'sd13, 8'sd16, 8'sd14, 8'sd23, 8'sd19, 8'sd47, 8'sd47, 8'sd20, 8'sd14, 8'sd10, 8'sd8, 8'sd1, 8'sd9, 8'sd24, 8'sd29, 8'sd18, -8'sd13, -8'sd14, 8'sd16, 8'sd63, 8'sd52, 8'sd25, 8'sd11, 8'sd9, 8'sd8, 8'sd16, 8'sd32, 8'sd36, 8'sd5, 8'sd4, -8'sd23, 8'sd11, 8'sd44, 8'sd51, 8'sd28, 8'sd18, 8'sd10, 8'sd13, 8'sd12, 8'sd24, 8'sd26, 8'sd8, 8'sd17, -8'sd3, 8'sd3, 8'sd29, 8'sd41, 8'sd32, 8'sd16, 8'sd10, 8'sd11, 8'sd8, 8'sd13, 8'sd16, 8'sd16, 8'sd9, 8'sd20, 8'sd10, 8'sd15, 8'sd28, 8'sd24, 8'sd8, 8'sd12, 8'sd16, 8'sd11, 8'sd8, 8'sd10, 8'sd18, 8'sd18, 8'sd9, 8'sd9, 8'sd19, 8'sd25, 8'sd29, 8'sd13, 8'sd8, -8'sd1, 8'sd15, 8'sd9, 8'sd10, 8'sd7, 8'sd19, 8'sd18, 8'sd19, 8'sd19, 8'sd11, 8'sd15, 8'sd5, 8'sd8, 8'sd4, 8'sd4, 8'sd14, 8'sd12, 8'sd9, 8'sd9, 8'sd20, 8'sd23, 8'sd20, 8'sd20, 8'sd26, 8'sd14, 8'sd12, 8'sd15, 8'sd21, 8'sd27, 8'sd13, 8'sd11, 8'sd11, 8'sd6, 8'sd8, 8'sd19, 8'sd12, 8'sd10, 8'sd18, 8'sd24, 8'sd9, 8'sd1, 8'sd22, 8'sd16, 8'sd13, 8'sd10, 8'sd9, 8'sd9, 8'sd5, 8'sd4, 8'sd5, 8'sd15, 8'sd15, 8'sd16, 8'sd14, 8'sd18, 8'sd16, 8'sd10, 8'sd8, 8'sd11, 8'sd8, 8'sd12, 8'sd8, 8'sd10, 8'sd11, 8'sd13, 8'sd12, 8'sd14, 8'sd11, 8'sd10, 8'sd10, 8'sd13, 8'sd10, 8'sd10,
    8'sd14, 8'sd15, 8'sd15, 8'sd11, 8'sd11, 8'sd14, 8'sd15, 8'sd15, 8'sd15, 8'sd11, 8'sd15, 8'sd14, 8'sd14, 8'sd12, 8'sd14, 8'sd11, 8'sd13, 8'sd19, 8'sd20, 8'sd23, 8'sd27, 8'sd24, 8'sd12, 8'sd15, 8'sd17, 8'sd15, 8'sd12, 8'sd12, 8'sd14, 8'sd9, 8'sd6, 8'sd14, 8'sd16, 8'sd20, 8'sd27, 8'sd20, 8'sd11, 8'sd13, 8'sd12, 8'sd18, 8'sd14, 8'sd12, 8'sd12, 8'sd11, -8'sd3, 8'sd9, 8'sd15, 8'sd7, 8'sd3, 8'sd23, 8'sd29, 8'sd5, 8'sd9, 8'sd14, 8'sd28, 8'sd12, 8'sd15, 8'sd10, -8'sd4, -8'sd2, 8'sd0, 8'sd11, 8'sd15, 8'sd21, 8'sd4, 8'sd6, 8'sd9, 8'sd36, 8'sd47, 8'sd12, 8'sd11, 8'sd11, 8'sd16, 8'sd32, 8'sd40, 8'sd41, 8'sd50, 8'sd13, -8'sd16, 8'sd3, 8'sd23, 8'sd38, 8'sd28, 8'sd15, 8'sd12, 8'sd13, 8'sd28, 8'sd46, 8'sd36, 8'sd26, 8'sd30, 8'sd26, 8'sd8, 8'sd9, 8'sd20, 8'sd25, 8'sd14, 8'sd14, 8'sd12, 8'sd10, 8'sd10, 8'sd7, 8'sd17, 8'sd14, 8'sd22, -8'sd1, 8'sd7, 8'sd1, 8'sd1, 8'sd22, 8'sd12, 8'sd12, 8'sd12, 8'sd6, 8'sd6, 8'sd11, 8'sd22, 8'sd26, 8'sd8, -8'sd3, 8'sd3, -8'sd1, 8'sd5, 8'sd16, 8'sd14, 8'sd14, 8'sd11, 8'sd9, 8'sd7, 8'sd13, 8'sd19, 8'sd39, 8'sd19, -8'sd2, 8'sd19, 8'sd20, 8'sd20, 8'sd22, 8'sd10, 8'sd14, 8'sd13, 8'sd8, 8'sd6, 8'sd6, 8'sd14, 8'sd23, 8'sd26, 8'sd2, 8'sd7, 8'sd7, 8'sd12, 8'sd23, 8'sd13, 8'sd11, 8'sd11, 8'sd10, 8'sd7, 8'sd5, 8'sd17, 8'sd27, 8'sd34, 8'sd11, 8'sd6, 8'sd0, 8'sd11, 8'sd13, 8'sd9, 8'sd13, 8'sd10, 8'sd13, 8'sd7, 8'sd9, 8'sd20, 8'sd25, 8'sd29, 8'sd18, 8'sd22, 8'sd18, 8'sd13, 8'sd10, 8'sd11, 8'sd15, 8'sd11, 8'sd14, 8'sd12, 8'sd11, 8'sd13, 8'sd17, 8'sd21, 8'sd17, 8'sd15, 8'sd13, 8'sd13, 8'sd13, 8'sd12, 8'sd14,
    8'sd19, 8'sd19, 8'sd19, 8'sd14, 8'sd16, 8'sd18, 8'sd18, 8'sd17, 8'sd17, 8'sd17, 8'sd17, 8'sd16, 8'sd16, 8'sd18, 8'sd19, 8'sd16, 8'sd18, 8'sd18, 8'sd17, 8'sd17, 8'sd19, 8'sd16, 8'sd15, 8'sd18, 8'sd13, 8'sd13, 8'sd16, 8'sd15, 8'sd16, 8'sd17, 8'sd17, 8'sd15, 8'sd10, 8'sd12, 8'sd19, 8'sd24, 8'sd36, 8'sd22, 8'sd18, 8'sd4, 8'sd19, 8'sd20, 8'sd16, 8'sd18, 8'sd17, 8'sd9, 8'sd4, 8'sd14, 8'sd6, 8'sd12, 8'sd30, 8'sd29, 8'sd22, 8'sd14, 8'sd7, 8'sd14, 8'sd17, 8'sd16, 8'sd17, 8'sd20, 8'sd22, 8'sd15, 8'sd18, -8'sd1, 8'sd10, 8'sd53, 8'sd24, 8'sd26, -8'sd13, 8'sd12, 8'sd16, 8'sd11, 8'sd14, 8'sd15, 8'sd23, 8'sd10, 8'sd7, -8'sd40, 8'sd42, 8'sd47, 8'sd30, 8'sd31, -8'sd13, 8'sd10, 8'sd15, 8'sd15, 8'sd8, 8'sd11, 8'sd8, -8'sd2, 8'sd1, 8'sd7, 8'sd38, 8'sd36, 8'sd39, 8'sd65, 8'sd50, 8'sd14, 8'sd18, 8'sd14, 8'sd21, 8'sd29, 8'sd2, 8'sd8, 8'sd15, 8'sd21, 8'sd20, 8'sd18, 8'sd9, 8'sd15, 8'sd26, 8'sd16, 8'sd16, 8'sd15, 8'sd15, 8'sd22, 8'sd29, 8'sd10, 8'sd23, 8'sd13, 8'sd24, 8'sd8, 8'sd11, 8'sd10, 8'sd11, 8'sd18, 8'sd18, 8'sd17, 8'sd4, 8'sd4, 8'sd20, 8'sd20, 8'sd12, 8'sd9, 8'sd8, 8'sd7, 8'sd0, -8'sd2, 8'sd14, 8'sd18, 8'sd15, 8'sd18, 8'sd13, 8'sd28, 8'sd13, 8'sd17, 8'sd18, 8'sd19, 8'sd4, 8'sd6, 8'sd2, -8'sd1, 8'sd14, 8'sd15, 8'sd18, 8'sd18, 8'sd8, 8'sd21, 8'sd8, 8'sd12, 8'sd22, 8'sd14, 8'sd4, 8'sd11, 8'sd11, 8'sd14, 8'sd20, 8'sd16, 8'sd18, 8'sd15, 8'sd13, 8'sd11, 8'sd9, 8'sd17, 8'sd17, 8'sd19, 8'sd16, 8'sd17, 8'sd12, 8'sd15, 8'sd16, 8'sd15, 8'sd17, 8'sd17, 8'sd14, 8'sd18, 8'sd17, 8'sd16, 8'sd14, 8'sd11, 8'sd14, 8'sd16, 8'sd16, 8'sd15, 8'sd15, 8'sd16,
    8'sd17, 8'sd14, 8'sd14, 8'sd14, 8'sd13, 8'sd16, 8'sd15, 8'sd15, 8'sd17, 8'sd15, 8'sd17, 8'sd15, 8'sd15, 8'sd16, 8'sd16, 8'sd15, 8'sd15, 8'sd12, 8'sd11, 8'sd10, 8'sd11, 8'sd11, 8'sd9, 8'sd14, 8'sd18, 8'sd17, 8'sd13, 8'sd13, 8'sd16, 8'sd13, 8'sd10, 8'sd0, 8'sd2, 8'sd9, 8'sd9, 8'sd6, 8'sd15, 8'sd16, 8'sd23, 8'sd34, 8'sd18, 8'sd17, 8'sd14, 8'sd13, 8'sd1, 8'sd6, 8'sd20, 8'sd27, 8'sd26, 8'sd8, 8'sd9, 8'sd16, 8'sd13, 8'sd25, 8'sd24, 8'sd14, 8'sd16, 8'sd12, 8'sd0, 8'sd11, 8'sd17, 8'sd32, 8'sd12, 8'sd14, 8'sd22, 8'sd21, 8'sd17, 8'sd14, 8'sd27, 8'sd15, 8'sd16, 8'sd13, 8'sd17, 8'sd24, 8'sd23, 8'sd46, 8'sd9, -8'sd15, 8'sd22, 8'sd4, 8'sd4, 8'sd5, 8'sd14, 8'sd15, 8'sd15, 8'sd17, 8'sd30, 8'sd44, 8'sd32, 8'sd33, -8'sd1, -8'sd12, 8'sd22, 8'sd28, 8'sd22, 8'sd22, 8'sd11, 8'sd13, 8'sd17, 8'sd16, 8'sd32, 8'sd35, 8'sd23, 8'sd17, -8'sd1, -8'sd24, 8'sd23, 8'sd13, 8'sd17, 8'sd23, 8'sd18, 8'sd13, 8'sd13, 8'sd10, 8'sd23, 8'sd22, 8'sd13, 8'sd12, -8'sd16, -8'sd3, 8'sd28, 8'sd18, 8'sd20, 8'sd2, 8'sd12, 8'sd13, 8'sd15, 8'sd7, 8'sd15, 8'sd15, 8'sd9, 8'sd0, -8'sd20, 8'sd21, 8'sd14, 8'sd14, 8'sd6, -8'sd2, 8'sd10, 8'sd12, 8'sd17, 8'sd12, 8'sd22, 8'sd15, -8'sd1, -8'sd4, 8'sd20, 8'sd19, 8'sd14, 8'sd10, 8'sd2, 8'sd16, 8'sd16, 8'sd15, 8'sd17, 8'sd11, 8'sd9, 8'sd4, 8'sd4, 8'sd5, 8'sd25, 8'sd19, 8'sd19, 8'sd17, 8'sd20, 8'sd20, 8'sd15, 8'sd13, 8'sd17, 8'sd12, 8'sd14, 8'sd8, 8'sd11, 8'sd13, 8'sd15, 8'sd17, 8'sd20, 8'sd20, 8'sd23, 8'sd17, 8'sd14, 8'sd17, 8'sd16, 8'sd13, 8'sd17, 8'sd17, 8'sd18, 8'sd21, 8'sd19, 8'sd19, 8'sd19, 8'sd19, 8'sd14, 8'sd18, 8'sd16, 8'sd17,
    8'sd13, 8'sd14, 8'sd12, 8'sd11, 8'sd10, 8'sd10, 8'sd12, 8'sd12, 8'sd12, 8'sd10, 8'sd14, 8'sd11, 8'sd10, 8'sd14, 8'sd12, 8'sd14, 8'sd12, 8'sd15, 8'sd13, 8'sd12, 8'sd18, 8'sd15, 8'sd12, 8'sd6, 8'sd8, 8'sd12, 8'sd10, 8'sd10, 8'sd13, 8'sd14, 8'sd13, 8'sd14, 8'sd18, 8'sd17, 8'sd9, 8'sd7, -8'sd9, 8'sd12, -8'sd1, -8'sd3, 8'sd12, 8'sd12, 8'sd11, 8'sd13, 8'sd10, 8'sd9, 8'sd18, 8'sd24, 8'sd45, 8'sd36, 8'sd37, 8'sd37, 8'sd37, -8'sd3, 8'sd3, 8'sd10, 8'sd13, 8'sd10, 8'sd1, 8'sd9, 8'sd21, 8'sd20, 8'sd35, 8'sd55, 8'sd42, 8'sd24, 8'sd16, 8'sd27, 8'sd14, 8'sd11, 8'sd13, 8'sd15, 8'sd12, 8'sd26, 8'sd23, 8'sd30, 8'sd41, 8'sd30, 8'sd22, 8'sd25, 8'sd27, 8'sd35, 8'sd24, 8'sd11, 8'sd12, 8'sd19, 8'sd31, 8'sd20, 8'sd21, 8'sd6, -8'sd22, 8'sd6, 8'sd14, 8'sd18, 8'sd16, 8'sd15, 8'sd5, 8'sd13, 8'sd14, 8'sd14, 8'sd17, 8'sd11, 8'sd2, 8'sd1, -8'sd11, -8'sd9, 8'sd4, -8'sd3, 8'sd13, -8'sd3, 8'sd4, 8'sd12, 8'sd12, 8'sd13, 8'sd12, -8'sd3, 8'sd3, 8'sd24, -8'sd4, -8'sd18, 8'sd1, 8'sd6, -8'sd6, -8'sd4, 8'sd5, 8'sd10, 8'sd14, 8'sd7, 8'sd12, 8'sd12, 8'sd18, 8'sd12, -8'sd4, 8'sd9, 8'sd9, 8'sd25, 8'sd22, 8'sd15, 8'sd7, 8'sd13, 8'sd10, 8'sd11, 8'sd19, 8'sd21, 8'sd20, -8'sd6, 8'sd2, 8'sd9, 8'sd8, 8'sd17, 8'sd21, 8'sd22, 8'sd14, 8'sd10, 8'sd13, 8'sd11, 8'sd15, 8'sd26, 8'sd30, 8'sd12, 8'sd8, 8'sd0, -8'sd4, -8'sd9, 8'sd3, 8'sd26, 8'sd14, 8'sd11, 8'sd11, 8'sd11, 8'sd17, 8'sd30, 8'sd34, 8'sd29, 8'sd31, 8'sd34, 8'sd38, 8'sd34, 8'sd21, 8'sd22, 8'sd15, 8'sd11, 8'sd13, 8'sd14, 8'sd15, 8'sd20, 8'sd24, 8'sd27, 8'sd32, 8'sd36, 8'sd33, 8'sd26, 8'sd16, 8'sd15, 8'sd12, 8'sd12,
    8'sd20, 8'sd16, 8'sd15, 8'sd19, 8'sd19, 8'sd17, 8'sd16, 8'sd19, 8'sd18, 8'sd16, 8'sd16, 8'sd17, 8'sd19, 8'sd17, 8'sd20, 8'sd20, 8'sd18, 8'sd16, 8'sd15, 8'sd12, 8'sd9, 8'sd9, 8'sd14, 8'sd21, 8'sd20, 8'sd23, 8'sd17, 8'sd17, 8'sd18, 8'sd18, 8'sd20, 8'sd19, 8'sd10, 8'sd2, 8'sd6, 8'sd16, 8'sd7, 8'sd13, 8'sd26, 8'sd27, 8'sd14, 8'sd18, 8'sd19, 8'sd18, 8'sd18, 8'sd17, 8'sd4, -8'sd1, -8'sd14, -8'sd25, -8'sd21, 8'sd2, 8'sd13, 8'sd20, 8'sd12, 8'sd14, 8'sd15, 8'sd16, 8'sd17, 8'sd3, -8'sd8, -8'sd19, -8'sd11, 8'sd0, 8'sd18, 8'sd4, 8'sd6, -8'sd8, -8'sd8, 8'sd11, 8'sd19, 8'sd18, 8'sd14, 8'sd17, 8'sd33, 8'sd54, 8'sd63, 8'sd26, 8'sd5, 8'sd6, 8'sd19, 8'sd2, -8'sd3, 8'sd15, 8'sd16, 8'sd16, 8'sd27, 8'sd39, 8'sd42, 8'sd26, 8'sd11, 8'sd17, 8'sd19, 8'sd13, 8'sd15, 8'sd27, 8'sd19, 8'sd14, 8'sd17, 8'sd16, 8'sd28, 8'sd22, 8'sd12, 8'sd7, 8'sd25, 8'sd22, 8'sd15, 8'sd18, 8'sd22, 8'sd26, 8'sd16, 8'sd15, 8'sd15, 8'sd12, -8'sd5, 8'sd14, 8'sd27, 8'sd23, 8'sd26, 8'sd17, 8'sd8, 8'sd18, 8'sd19, 8'sd4, -8'sd1, 8'sd15, 8'sd18, 8'sd13, -8'sd13, -8'sd22, 8'sd18, 8'sd23, 8'sd28, 8'sd15, 8'sd12, 8'sd18, 8'sd12, 8'sd0, 8'sd0, 8'sd17, 8'sd18, 8'sd12, 8'sd0, -8'sd3, 8'sd1, 8'sd10, 8'sd19, 8'sd24, 8'sd22, 8'sd20, 8'sd2, -8'sd1, 8'sd13, 8'sd19, 8'sd15, 8'sd17, 8'sd20, 8'sd20, 8'sd15, 8'sd15, 8'sd20, 8'sd25, 8'sd23, 8'sd24, 8'sd8, 8'sd6, 8'sd13, 8'sd17, 8'sd18, 8'sd16, 8'sd18, 8'sd15, 8'sd12, 8'sd20, 8'sd10, 8'sd9, 8'sd6, 8'sd9, 8'sd9, 8'sd14, 8'sd13, 8'sd16, 8'sd15, 8'sd18, 8'sd18, 8'sd17, 8'sd16, 8'sd15, 8'sd10, 8'sd5, 8'sd8, 8'sd12, 8'sd12, 8'sd17, 8'sd18, 8'sd15,
    8'sd19, 8'sd16, 8'sd16, 8'sd17, 8'sd16, 8'sd18, 8'sd16, 8'sd19, 8'sd15, 8'sd17, 8'sd18, 8'sd18, 8'sd19, 8'sd17, 8'sd18, 8'sd15, 8'sd17, 8'sd18, 8'sd17, 8'sd18, 8'sd21, 8'sd22, 8'sd26, 8'sd19, 8'sd18, 8'sd20, 8'sd17, 8'sd18, 8'sd20, 8'sd19, 8'sd20, 8'sd14, 8'sd15, 8'sd11, 8'sd9, 8'sd8, -8'sd2, 8'sd5, 8'sd16, 8'sd19, 8'sd10, 8'sd19, 8'sd16, 8'sd14, 8'sd9, -8'sd7, -8'sd11, -8'sd2, -8'sd4, 8'sd10, 8'sd5, 8'sd4, 8'sd9, 8'sd6, 8'sd6, 8'sd14, 8'sd16, 8'sd14, -8'sd6, -8'sd10, -8'sd11, 8'sd2, 8'sd16, 8'sd17, -8'sd5, 8'sd5, 8'sd8, -8'sd7, -8'sd2, 8'sd16, 8'sd19, 8'sd11, 8'sd10, 8'sd9, 8'sd11, 8'sd3, -8'sd11, 8'sd3, 8'sd11, 8'sd9, 8'sd7, -8'sd9, -8'sd1, 8'sd15, 8'sd18, 8'sd18, 8'sd30, 8'sd35, 8'sd26, 8'sd21, 8'sd48, 8'sd45, 8'sd17, 8'sd33, 8'sd37, 8'sd16, 8'sd12, 8'sd16, 8'sd17, 8'sd18, 8'sd34, 8'sd39, 8'sd32, 8'sd27, 8'sd36, 8'sd30, 8'sd25, 8'sd19, 8'sd21, 8'sd9, 8'sd18, 8'sd19, 8'sd19, 8'sd18, 8'sd26, 8'sd28, 8'sd9, 8'sd20, 8'sd27, 8'sd34, 8'sd23, 8'sd14, 8'sd13, 8'sd9, 8'sd14, 8'sd18, 8'sd19, 8'sd15, 8'sd5, 8'sd8, 8'sd28, 8'sd30, 8'sd36, 8'sd43, 8'sd27, 8'sd18, 8'sd11, 8'sd7, 8'sd21, 8'sd20, 8'sd16, 8'sd17, 8'sd2, -8'sd22, -8'sd17, 8'sd1, 8'sd8, 8'sd7, 8'sd6, 8'sd12, 8'sd0, 8'sd8, 8'sd18, 8'sd18, 8'sd18, 8'sd17, 8'sd12, 8'sd0, -8'sd9, -8'sd27, -8'sd28, -8'sd19, -8'sd17, -8'sd4, 8'sd6, 8'sd15, 8'sd19, 8'sd15, 8'sd18, 8'sd17, 8'sd15, 8'sd15, 8'sd15, 8'sd9, -8'sd1, -8'sd4, 8'sd16, 8'sd16, 8'sd30, 8'sd20, 8'sd19, 8'sd19, 8'sd18, 8'sd20, 8'sd17, 8'sd18, 8'sd13, 8'sd14, 8'sd20, 8'sd21, 8'sd16, 8'sd14, 8'sd19, 8'sd18, 8'sd17, 8'sd16,
    8'sd12, 8'sd13, 8'sd13, 8'sd13, 8'sd11, 8'sd11, 8'sd14, 8'sd12, 8'sd10, 8'sd11, 8'sd12, 8'sd11, 8'sd15, 8'sd15, 8'sd13, 8'sd15, 8'sd14, 8'sd13, 8'sd15, 8'sd22, 8'sd26, 8'sd19, 8'sd15, 8'sd17, 8'sd15, 8'sd14, 8'sd13, 8'sd13, 8'sd14, 8'sd12, 8'sd15, 8'sd20, 8'sd24, 8'sd30, 8'sd24, 8'sd2, 8'sd15, 8'sd23, 8'sd21, 8'sd15, 8'sd19, 8'sd13, 8'sd14, 8'sd11, 8'sd16, 8'sd18, 8'sd31, 8'sd12, 8'sd12, 8'sd23, 8'sd18, 8'sd4, 8'sd7, 8'sd13, 8'sd19, 8'sd11, 8'sd12, 8'sd10, 8'sd5, 8'sd10, 8'sd15, 8'sd16, 8'sd7, 8'sd0, -8'sd1, 8'sd1, 8'sd4, 8'sd7, 8'sd6, 8'sd15, 8'sd11, 8'sd7, 8'sd8, 8'sd20, 8'sd34, 8'sd20, -8'sd16, -8'sd18, 8'sd1, 8'sd4, 8'sd2, -8'sd3, 8'sd2, 8'sd14, 8'sd11, 8'sd10, 8'sd6, 8'sd4, 8'sd20, 8'sd43, 8'sd26, 8'sd12, 8'sd18, 8'sd20, 8'sd16, 8'sd8, 8'sd15, 8'sd15, 8'sd15, 8'sd15, 8'sd6, 8'sd15, 8'sd16, 8'sd30, 8'sd34, 8'sd19, 8'sd25, 8'sd11, 8'sd9, 8'sd12, 8'sd14, 8'sd14, 8'sd12, 8'sd14, 8'sd12, 8'sd6, 8'sd19, 8'sd26, 8'sd43, 8'sd22, 8'sd27, 8'sd29, 8'sd24, 8'sd24, 8'sd22, 8'sd16, 8'sd15, 8'sd19, 8'sd27, 8'sd19, -8'sd1, 8'sd12, 8'sd15, 8'sd11, 8'sd17, 8'sd16, 8'sd24, 8'sd23, 8'sd24, 8'sd14, 8'sd11, 8'sd19, 8'sd24, 8'sd13, 8'sd10, -8'sd3, 8'sd20, 8'sd28, 8'sd17, 8'sd25, 8'sd24, 8'sd31, 8'sd15, 8'sd15, 8'sd13, 8'sd17, 8'sd22, 8'sd12, 8'sd22, 8'sd18, 8'sd8, 8'sd13, 8'sd21, 8'sd41, 8'sd35, 8'sd23, 8'sd16, 8'sd13, 8'sd12, 8'sd15, 8'sd13, 8'sd9, 8'sd12, 8'sd19, 8'sd18, 8'sd20, 8'sd14, 8'sd20, 8'sd21, 8'sd19, 8'sd15, 8'sd14, 8'sd12, 8'sd11, 8'sd14, 8'sd13, 8'sd14, 8'sd13, 8'sd12, 8'sd13, 8'sd6, 8'sd5, 8'sd13, 8'sd14, 8'sd15, 8'sd12,
    8'sd13, 8'sd14, 8'sd12, 8'sd13, 8'sd13, 8'sd17, 8'sd13, 8'sd14, 8'sd16, 8'sd14, 8'sd16, 8'sd13, 8'sd14, 8'sd14, 8'sd13, 8'sd16, 8'sd14, 8'sd12, 8'sd17, 8'sd14, 8'sd7, 8'sd10, 8'sd9, 8'sd15, 8'sd18, 8'sd17, 8'sd14, 8'sd16, 8'sd14, 8'sd15, 8'sd13, 8'sd13, 8'sd13, 8'sd12, -8'sd1, -8'sd4, 8'sd1, 8'sd3, 8'sd20, 8'sd30, 8'sd20, 8'sd17, 8'sd15, 8'sd13, 8'sd11, 8'sd19, 8'sd26, 8'sd32, 8'sd20, -8'sd1, -8'sd13, 8'sd5, 8'sd9, 8'sd29, 8'sd35, 8'sd16, 8'sd15, 8'sd13, 8'sd15, 8'sd13, 8'sd17, 8'sd22, 8'sd46, 8'sd0, -8'sd28, -8'sd12, 8'sd6, 8'sd10, 8'sd38, 8'sd15, 8'sd15, 8'sd14, 8'sd14, 8'sd20, 8'sd21, 8'sd18, 8'sd34, 8'sd42, 8'sd1, -8'sd18, -8'sd8, 8'sd3, 8'sd22, 8'sd18, 8'sd12, 8'sd12, 8'sd15, 8'sd24, 8'sd17, 8'sd14, 8'sd35, 8'sd33, 8'sd18, 8'sd10, 8'sd13, 8'sd6, 8'sd12, 8'sd13, 8'sd14, 8'sd14, 8'sd8, 8'sd7, 8'sd14, 8'sd28, 8'sd28, 8'sd37, 8'sd4, 8'sd12, 8'sd9, 8'sd8, 8'sd16, 8'sd14, 8'sd13, 8'sd12, 8'sd2, 8'sd10, 8'sd19, 8'sd21, 8'sd37, 8'sd27, 8'sd13, 8'sd9, 8'sd16, 8'sd17, 8'sd19, 8'sd13, 8'sd16, 8'sd13, 8'sd15, 8'sd17, 8'sd24, 8'sd20, 8'sd14, 8'sd18, 8'sd14, 8'sd14, 8'sd20, 8'sd24, 8'sd13, 8'sd16, 8'sd17, 8'sd9, 8'sd8, 8'sd19, 8'sd20, 8'sd11, 8'sd4, 8'sd21, 8'sd20, 8'sd20, 8'sd18, 8'sd17, 8'sd11, 8'sd12, 8'sd17, 8'sd11, 8'sd12, 8'sd20, 8'sd17, 8'sd10, 8'sd14, 8'sd9, 8'sd23, 8'sd16, 8'sd15, 8'sd13, 8'sd12, 8'sd16, 8'sd16, 8'sd14, 8'sd5, -8'sd1, 8'sd5, 8'sd8, 8'sd9, 8'sd14, 8'sd19, 8'sd26, 8'sd12, 8'sd16, 8'sd16, 8'sd14, 8'sd15, 8'sd14, 8'sd12, 8'sd12, 8'sd10, 8'sd7, 8'sd1, 8'sd3, 8'sd9, 8'sd10, 8'sd15, 8'sd14, 8'sd13, 8'sd13,
    8'sd14, 8'sd16, 8'sd14, 8'sd14, 8'sd17, 8'sd16, 8'sd16, 8'sd13, 8'sd16, 8'sd17, 8'sd14, 8'sd13, 8'sd15, 8'sd14, 8'sd16, 8'sd17, 8'sd17, 8'sd14, 8'sd12, 8'sd13, 8'sd11, 8'sd15, 8'sd12, 8'sd13, 8'sd16, 8'sd15, 8'sd17, 8'sd16, 8'sd12, 8'sd15, 8'sd18, 8'sd17, 8'sd9, 8'sd2, 8'sd1, 8'sd18, 8'sd7, 8'sd9, 8'sd4, 8'sd11, 8'sd13, 8'sd13, 8'sd17, 8'sd19, 8'sd29, 8'sd27, 8'sd24, 8'sd25, 8'sd13, 8'sd27, 8'sd19, 8'sd19, 8'sd21, 8'sd7, 8'sd7, 8'sd14, 8'sd14, 8'sd20, 8'sd29, 8'sd25, 8'sd23, 8'sd24, 8'sd6, 8'sd43, 8'sd17, 8'sd28, 8'sd21, 8'sd13, 8'sd7, 8'sd12, 8'sd18, 8'sd29, 8'sd19, 8'sd1, 8'sd3, 8'sd11, 8'sd6, 8'sd63, 8'sd55, 8'sd38, 8'sd29, 8'sd12, 8'sd14, 8'sd17, 8'sd15, 8'sd21, 8'sd4, 8'sd3, -8'sd2, -8'sd10, -8'sd18, 8'sd5, 8'sd11, 8'sd9, 8'sd12, 8'sd19, 8'sd17, 8'sd15, 8'sd15, 8'sd14, 8'sd9, 8'sd0, 8'sd4, -8'sd2, -8'sd4, -8'sd3, 8'sd0, 8'sd19, 8'sd33, 8'sd33, 8'sd15, 8'sd15, 8'sd12, 8'sd17, 8'sd13, 8'sd3, 8'sd11, 8'sd0, -8'sd6, 8'sd6, 8'sd10, 8'sd17, 8'sd25, 8'sd23, 8'sd14, 8'sd14, 8'sd17, 8'sd22, 8'sd15, 8'sd1, 8'sd12, 8'sd7, 8'sd3, 8'sd12, 8'sd10, 8'sd12, 8'sd9, 8'sd11, 8'sd12, 8'sd13, 8'sd12, 8'sd20, 8'sd23, 8'sd25, 8'sd30, 8'sd24, 8'sd35, 8'sd24, 8'sd12, 8'sd0, 8'sd1, -8'sd1, 8'sd13, 8'sd17, 8'sd13, 8'sd16, 8'sd26, 8'sd37, 8'sd20, 8'sd14, 8'sd14, 8'sd24, 8'sd20, 8'sd16, -8'sd2, 8'sd3, 8'sd11, 8'sd13, 8'sd12, 8'sd14, 8'sd18, 8'sd24, 8'sd20, 8'sd18, 8'sd16, 8'sd6, 8'sd11, 8'sd7, 8'sd1, 8'sd8, 8'sd16, 8'sd14, 8'sd14, 8'sd17, 8'sd12, 8'sd12, 8'sd14, 8'sd12, 8'sd13, 8'sd22, 8'sd20, 8'sd22, 8'sd14, 8'sd16, 8'sd16, 8'sd14,
    8'sd19, 8'sd16, 8'sd17, 8'sd15, 8'sd16, 8'sd16, 8'sd14, 8'sd16, 8'sd17, 8'sd15, 8'sd15, 8'sd19, 8'sd16, 8'sd15, 8'sd16, 8'sd16, 8'sd15, 8'sd18, 8'sd20, 8'sd20, 8'sd17, 8'sd9, 8'sd10, 8'sd8, 8'sd14, 8'sd17, 8'sd16, 8'sd19, 8'sd19, 8'sd17, 8'sd15, 8'sd14, 8'sd17, 8'sd15, 8'sd14, 8'sd13, 8'sd4, 8'sd7, 8'sd14, 8'sd12, 8'sd19, 8'sd18, 8'sd18, 8'sd14, 8'sd18, 8'sd18, 8'sd21, 8'sd27, 8'sd19, 8'sd12, 8'sd6, 8'sd19, 8'sd16, 8'sd14, 8'sd21, 8'sd19, 8'sd17, 8'sd18, 8'sd17, 8'sd16, 8'sd23, 8'sd32, 8'sd31, 8'sd32, 8'sd21, 8'sd21, 8'sd18, 8'sd18, 8'sd21, 8'sd18, 8'sd16, 8'sd17, 8'sd10, 8'sd15, 8'sd18, 8'sd12, 8'sd19, 8'sd15, 8'sd8, 8'sd5, -8'sd4, -8'sd2, 8'sd19, 8'sd20, 8'sd19, 8'sd15, -8'sd3, -8'sd15, -8'sd18, -8'sd28, -8'sd30, -8'sd11, -8'sd6, -8'sd9, -8'sd4, 8'sd0, 8'sd14, 8'sd18, 8'sd15, 8'sd16, -8'sd9, -8'sd31, -8'sd10, 8'sd3, 8'sd17, 8'sd10, 8'sd5, 8'sd7, 8'sd16, 8'sd7, 8'sd19, 8'sd25, 8'sd19, 8'sd11, 8'sd2, 8'sd16, 8'sd26, 8'sd19, 8'sd25, 8'sd21, 8'sd11, 8'sd3, 8'sd20, 8'sd14, 8'sd26, 8'sd24, 8'sd19, 8'sd13, 8'sd16, 8'sd20, 8'sd27, 8'sd21, 8'sd24, 8'sd27, 8'sd15, 8'sd7, 8'sd2, 8'sd8, 8'sd28, 8'sd21, 8'sd15, 8'sd17, 8'sd16, 8'sd12, 8'sd18, 8'sd20, 8'sd21, 8'sd22, 8'sd14, 8'sd15, 8'sd4, 8'sd20, 8'sd26, 8'sd19, 8'sd18, 8'sd15, 8'sd12, 8'sd18, 8'sd18, 8'sd18, 8'sd18, 8'sd20, 8'sd10, 8'sd17, 8'sd23, 8'sd27, 8'sd19, 8'sd16, 8'sd19, 8'sd15, 8'sd12, 8'sd8, 8'sd9, 8'sd12, 8'sd8, 8'sd12, 8'sd17, 8'sd20, 8'sd17, 8'sd17, 8'sd17, 8'sd17, 8'sd15, 8'sd18, 8'sd19, 8'sd17, 8'sd17, 8'sd22, 8'sd16, 8'sd22, 8'sd19, 8'sd16, 8'sd16, 8'sd16, 8'sd19, 8'sd15,
    8'sd16, 8'sd15, 8'sd18, 8'sd17, 8'sd18, 8'sd15, 8'sd17, 8'sd14, 8'sd17, 8'sd15, 8'sd17, 8'sd17, 8'sd14, 8'sd17, 8'sd15, 8'sd17, 8'sd15, 8'sd17, 8'sd15, 8'sd16, 8'sd15, 8'sd15, 8'sd14, 8'sd13, 8'sd14, 8'sd15, 8'sd17, 8'sd16, 8'sd17, 8'sd15, 8'sd16, 8'sd20, 8'sd19, 8'sd6, -8'sd4, -8'sd12, -8'sd15, -8'sd7, 8'sd3, 8'sd11, 8'sd17, 8'sd16, 8'sd14, 8'sd20, 8'sd24, 8'sd21, 8'sd27, 8'sd17, 8'sd31, 8'sd17, 8'sd20, 8'sd12, 8'sd13, 8'sd5, 8'sd12, 8'sd17, 8'sd16, 8'sd19, 8'sd20, 8'sd18, 8'sd20, 8'sd25, 8'sd27, 8'sd21, 8'sd18, 8'sd24, 8'sd17, 8'sd24, 8'sd10, 8'sd17, 8'sd15, 8'sd25, 8'sd17, 8'sd15, 8'sd18, 8'sd20, 8'sd15, 8'sd20, 8'sd21, 8'sd29, 8'sd35, 8'sd17, 8'sd9, 8'sd17, 8'sd19, 8'sd20, 8'sd16, 8'sd17, 8'sd5, 8'sd11, 8'sd13, 8'sd38, 8'sd32, 8'sd19, 8'sd13, 8'sd10, 8'sd10, 8'sd18, 8'sd15, 8'sd19, 8'sd9, 8'sd7, 8'sd10, 8'sd10, 8'sd14, 8'sd23, 8'sd22, 8'sd27, 8'sd21, 8'sd11, 8'sd16, 8'sd17, 8'sd16, 8'sd20, 8'sd17, 8'sd12, 8'sd16, 8'sd9, 8'sd8, 8'sd10, 8'sd20, 8'sd17, 8'sd24, 8'sd19, 8'sd14, 8'sd15, 8'sd18, 8'sd17, 8'sd13, -8'sd13, -8'sd10, -8'sd6, -8'sd8, 8'sd2, 8'sd4, 8'sd6, 8'sd16, 8'sd8, 8'sd11, 8'sd14, 8'sd17, 8'sd19, 8'sd5, -8'sd13, -8'sd7, -8'sd6, -8'sd5, -8'sd3, -8'sd1, 8'sd4, 8'sd8, -8'sd2, 8'sd12, 8'sd18, 8'sd18, 8'sd19, 8'sd20, 8'sd18, 8'sd8, 8'sd7, -8'sd3, 8'sd2, -8'sd4, -8'sd10, -8'sd6, 8'sd2, 8'sd13, 8'sd14, 8'sd16, 8'sd17, 8'sd31, 8'sd37, 8'sd23, 8'sd26, 8'sd24, 8'sd16, 8'sd16, 8'sd4, 8'sd13, 8'sd16, 8'sd14, 8'sd16, 8'sd14, 8'sd17, 8'sd18, 8'sd15, 8'sd18, 8'sd18, 8'sd20, 8'sd24, 8'sd24, 8'sd22, 8'sd18, 8'sd18, 8'sd14, 8'sd17,
    8'sd10, 8'sd12, 8'sd13, 8'sd8, 8'sd10, 8'sd9, 8'sd11, 8'sd11, 8'sd10, 8'sd13, 8'sd12, 8'sd10, 8'sd12, 8'sd12, 8'sd10, 8'sd8, 8'sd11, 8'sd8, 8'sd15, 8'sd21, 8'sd26, 8'sd19, 8'sd23, 8'sd17, 8'sd10, 8'sd14, 8'sd11, 8'sd12, 8'sd9, 8'sd10, 8'sd7, 8'sd7, 8'sd19, 8'sd17, 8'sd7, 8'sd4, 8'sd9, 8'sd3, 8'sd9, 8'sd15, 8'sd12, 8'sd12, 8'sd12, 8'sd10, 8'sd5, 8'sd16, 8'sd14, 8'sd8, 8'sd15, 8'sd9, 8'sd9, 8'sd13, 8'sd4, 8'sd9, 8'sd7, 8'sd9, 8'sd10, 8'sd13, 8'sd13, 8'sd17, 8'sd9, 8'sd17, 8'sd25, 8'sd26, 8'sd26, 8'sd13, 8'sd12, 8'sd9, -8'sd3, 8'sd9, 8'sd12, 8'sd17, 8'sd31, 8'sd25, 8'sd9, 8'sd11, -8'sd1, -8'sd6, 8'sd11, 8'sd12, 8'sd19, 8'sd25, 8'sd13, 8'sd12, 8'sd9, 8'sd20, 8'sd36, 8'sd32, 8'sd8, 8'sd8, -8'sd6, -8'sd20, -8'sd2, 8'sd5, 8'sd31, 8'sd46, 8'sd28, 8'sd9, 8'sd13, 8'sd13, 8'sd31, 8'sd55, 8'sd44, 8'sd18, -8'sd17, 8'sd1, 8'sd29, 8'sd34, 8'sd27, 8'sd23, 8'sd19, 8'sd10, 8'sd10, 8'sd10, 8'sd19, 8'sd34, 8'sd63, 8'sd58, 8'sd15, 8'sd28, 8'sd29, 8'sd18, 8'sd14, 8'sd5, 8'sd18, 8'sd13, 8'sd12, 8'sd3, 8'sd5, -8'sd1, 8'sd7, 8'sd41, 8'sd50, 8'sd23, 8'sd8, 8'sd18, 8'sd6, 8'sd13, 8'sd22, 8'sd11, 8'sd10, 8'sd9, 8'sd7, 8'sd6, 8'sd2, 8'sd10, 8'sd20, 8'sd25, 8'sd18, 8'sd10, 8'sd13, 8'sd29, 8'sd20, 8'sd10, 8'sd10, 8'sd11, 8'sd7, 8'sd15, 8'sd18, 8'sd13, 8'sd11, 8'sd6, 8'sd5, 8'sd21, 8'sd26, 8'sd27, 8'sd16, 8'sd12, 8'sd9, 8'sd11, 8'sd11, 8'sd6, 8'sd3, 8'sd7, 8'sd11, 8'sd18, 8'sd16, 8'sd15, 8'sd16, 8'sd12, 8'sd9, 8'sd12, 8'sd10, 8'sd10, 8'sd9, 8'sd11, 8'sd10, 8'sd13, 8'sd19, 8'sd18, 8'sd13, 8'sd15, 8'sd13, 8'sd12, 8'sd8, 8'sd12,
    8'sd13, 8'sd14, 8'sd16, 8'sd14, 8'sd16, 8'sd16, 8'sd15, 8'sd18, 8'sd15, 8'sd14, 8'sd17, 8'sd15, 8'sd14, 8'sd14, 8'sd16, 8'sd15, 8'sd15, 8'sd14, 8'sd4, -8'sd1, 8'sd1, 8'sd4, 8'sd3, 8'sd7, 8'sd7, 8'sd10, 8'sd14, 8'sd16, 8'sd14, 8'sd18, 8'sd19, 8'sd20, 8'sd13, 8'sd14, 8'sd23, 8'sd22, 8'sd12, 8'sd10, 8'sd9, 8'sd12, 8'sd17, 8'sd15, 8'sd16, 8'sd15, 8'sd22, 8'sd16, 8'sd21, 8'sd20, 8'sd14, 8'sd8, 8'sd4, -8'sd2, 8'sd9, 8'sd21, 8'sd17, 8'sd14, 8'sd17, 8'sd14, 8'sd24, 8'sd23, 8'sd15, 8'sd12, 8'sd14, 8'sd12, 8'sd16, 8'sd32, 8'sd25, 8'sd36, 8'sd27, 8'sd17, 8'sd14, 8'sd17, 8'sd17, 8'sd17, 8'sd16, 8'sd28, 8'sd28, 8'sd48, 8'sd37, 8'sd26, 8'sd27, 8'sd20, 8'sd24, 8'sd16, 8'sd15, 8'sd16, 8'sd15, 8'sd12, 8'sd23, 8'sd21, 8'sd28, 8'sd30, 8'sd26, 8'sd19, 8'sd19, 8'sd0, 8'sd16, 8'sd20, 8'sd17, 8'sd17, 8'sd12, -8'sd8, 8'sd11, 8'sd17, 8'sd21, 8'sd31, 8'sd40, 8'sd19, 8'sd3, 8'sd6, 8'sd9, 8'sd16, 8'sd15, 8'sd24, 8'sd20, 8'sd4, 8'sd2, -8'sd4, 8'sd33, 8'sd45, 8'sd16, -8'sd6, 8'sd5, 8'sd21, 8'sd14, 8'sd14, 8'sd14, 8'sd24, 8'sd24, 8'sd17, 8'sd6, 8'sd2, 8'sd6, -8'sd7, -8'sd18, -8'sd2, 8'sd1, 8'sd8, 8'sd8, 8'sd13, 8'sd13, 8'sd18, 8'sd13, 8'sd16, 8'sd7, 8'sd6, 8'sd0, 8'sd3, 8'sd9, 8'sd6, 8'sd2, 8'sd2, 8'sd8, 8'sd14, 8'sd18, 8'sd18, 8'sd12, 8'sd16, 8'sd10, 8'sd6, 8'sd15, 8'sd19, 8'sd20, 8'sd28, 8'sd21, 8'sd18, 8'sd15, 8'sd16, 8'sd15, 8'sd18, 8'sd17, 8'sd17, 8'sd21, 8'sd22, 8'sd6, 8'sd15, 8'sd14, 8'sd17, 8'sd17, 8'sd17, 8'sd15, 8'sd13, 8'sd13, 8'sd17, 8'sd13, 8'sd14, 8'sd17, 8'sd16, 8'sd19, 8'sd12, 8'sd15, 8'sd12, 8'sd15, 8'sd17, 8'sd17, 8'sd13,
    8'sd19, 8'sd22, 8'sd21, 8'sd18, 8'sd21, 8'sd21, 8'sd19, 8'sd20, 8'sd18, 8'sd18, 8'sd19, 8'sd19, 8'sd20, 8'sd21, 8'sd22, 8'sd20, 8'sd21, 8'sd21, 8'sd17, 8'sd8, 8'sd5, 8'sd9, 8'sd10, 8'sd15, 8'sd19, 8'sd21, 8'sd18, 8'sd21, 8'sd20, 8'sd19, 8'sd19, 8'sd16, 8'sd1, -8'sd6, -8'sd3, 8'sd6, 8'sd3, 8'sd9, 8'sd18, 8'sd26, 8'sd15, 8'sd20, 8'sd19, 8'sd20, 8'sd18, 8'sd3, -8'sd9, 8'sd1, 8'sd14, 8'sd6, 8'sd8, 8'sd16, 8'sd11, 8'sd19, 8'sd21, 8'sd20, 8'sd21, 8'sd17, 8'sd14, 8'sd3, -8'sd2, -8'sd1, 8'sd22, 8'sd27, 8'sd23, 8'sd17, 8'sd16, 8'sd15, 8'sd37, 8'sd21, 8'sd18, 8'sd19, 8'sd14, 8'sd7, 8'sd7, 8'sd10, 8'sd24, 8'sd33, 8'sd11, 8'sd0, 8'sd12, 8'sd30, 8'sd45, 8'sd23, 8'sd19, 8'sd19, 8'sd22, 8'sd19, 8'sd12, 8'sd11, 8'sd24, 8'sd20, 8'sd6, -8'sd32, -8'sd35, -8'sd20, 8'sd8, 8'sd22, 8'sd21, 8'sd22, 8'sd19, 8'sd13, 8'sd18, 8'sd14, 8'sd12, 8'sd13, 8'sd16, 8'sd13, -8'sd12, -8'sd8, 8'sd13, 8'sd17, 8'sd21, 8'sd17, 8'sd18, 8'sd11, 8'sd4, 8'sd9, 8'sd13, 8'sd23, 8'sd13, 8'sd15, -8'sd7, 8'sd0, 8'sd9, 8'sd19, 8'sd22, 8'sd17, 8'sd19, 8'sd21, 8'sd7, 8'sd8, 8'sd23, 8'sd15, 8'sd12, 8'sd16, -8'sd1, 8'sd3, 8'sd13, 8'sd20, 8'sd21, 8'sd14, 8'sd4, 8'sd8, 8'sd18, 8'sd15, 8'sd9, 8'sd15, 8'sd17, 8'sd17, 8'sd4, 8'sd10, 8'sd19, 8'sd22, 8'sd21, 8'sd19, 8'sd19, 8'sd9, 8'sd19, 8'sd15, 8'sd9, 8'sd7, 8'sd21, 8'sd24, 8'sd12, 8'sd17, 8'sd18, 8'sd21, 8'sd20, 8'sd19, 8'sd14, 8'sd11, 8'sd8, 8'sd12, 8'sd10, 8'sd5, 8'sd8, 8'sd17, 8'sd16, 8'sd19, 8'sd19, 8'sd18, 8'sd20, 8'sd18, 8'sd21, 8'sd16, 8'sd14, 8'sd16, 8'sd15, 8'sd15, 8'sd12, 8'sd17, 8'sd17, 8'sd22, 8'sd22, 8'sd20,
    8'sd13, 8'sd11, 8'sd13, 8'sd15, 8'sd11, 8'sd15, 8'sd12, 8'sd13, 8'sd15, 8'sd13, 8'sd11, 8'sd11, 8'sd12, 8'sd11, 8'sd10, 8'sd10, 8'sd15, 8'sd14, 8'sd19, 8'sd27, 8'sd31, 8'sd31, 8'sd26, 8'sd19, 8'sd13, 8'sd13, 8'sd13, 8'sd10, 8'sd14, 8'sd13, 8'sd13, 8'sd20, 8'sd28, 8'sd27, 8'sd24, 8'sd23, 8'sd22, 8'sd13, 8'sd6, 8'sd7, 8'sd14, 8'sd15, 8'sd12, 8'sd12, 8'sd10, 8'sd16, 8'sd23, 8'sd11, 8'sd14, 8'sd9, 8'sd5, 8'sd8, 8'sd5, 8'sd8, 8'sd17, 8'sd14, 8'sd14, 8'sd9, 8'sd3, 8'sd17, 8'sd20, 8'sd11, 8'sd3, 8'sd17, 8'sd9, 8'sd7, 8'sd18, 8'sd16, 8'sd24, 8'sd13, 8'sd11, 8'sd8, 8'sd11, 8'sd17, 8'sd4, 8'sd12, 8'sd23, 8'sd12, 8'sd7, 8'sd0, 8'sd9, 8'sd10, 8'sd22, 8'sd12, 8'sd14, 8'sd11, 8'sd2, -8'sd9, -8'sd1, 8'sd24, 8'sd18, -8'sd1, 8'sd2, 8'sd7, 8'sd7, 8'sd16, 8'sd22, 8'sd11, 8'sd12, 8'sd12, 8'sd9, 8'sd8, 8'sd14, 8'sd18, 8'sd11, 8'sd14, 8'sd3, 8'sd14, 8'sd18, 8'sd26, 8'sd33, 8'sd14, 8'sd14, 8'sd17, 8'sd26, 8'sd23, 8'sd3, 8'sd9, -8'sd3, 8'sd6, 8'sd10, 8'sd19, 8'sd14, 8'sd42, 8'sd38, 8'sd14, 8'sd12, 8'sd14, 8'sd26, 8'sd41, 8'sd40, 8'sd42, 8'sd19, 8'sd12, 8'sd20, 8'sd22, 8'sd17, 8'sd44, 8'sd29, 8'sd14, 8'sd11, 8'sd16, 8'sd26, 8'sd26, 8'sd40, 8'sd47, 8'sd34, 8'sd22, 8'sd18, 8'sd24, 8'sd20, 8'sd28, 8'sd18, 8'sd14, 8'sd14, 8'sd16, 8'sd10, 8'sd1, 8'sd9, 8'sd16, 8'sd26, 8'sd22, 8'sd19, 8'sd19, 8'sd25, 8'sd16, 8'sd15, 8'sd12, 8'sd14, 8'sd13, 8'sd7, 8'sd3, 8'sd0, 8'sd2, 8'sd2, 8'sd10, 8'sd11, 8'sd11, 8'sd5, 8'sd12, 8'sd12, 8'sd11, 8'sd10, 8'sd10, 8'sd11, 8'sd13, 8'sd10, 8'sd9, 8'sd10, 8'sd8, 8'sd9, 8'sd12, 8'sd9, 8'sd12, 8'sd10, 8'sd12
    };

    localparam signed [8*30-1:0] biases_HL_param = {
    8'sd20, 8'sd19, 8'sd16, 8'sd10, 8'sd18, 8'sd3, 8'sd2, 8'sd8, 8'sd17, 8'sd13, 8'sd14, 8'sd12, 8'sd18, 8'sd4, 8'sd24, 8'sd20, 8'sd10, 8'sd15, 8'sd20, 8'sd5, 8'sd7, 8'sd18, 8'sd14, 8'sd15, 8'sd9, 8'sd9, 8'sd23, 8'sd11, 8'sd0, 8'sd18
    };


    // Assign values to weights and biases
    always @(*) begin
        integer i, j;

        // Assign weights from the flattened localparam to the output
        for (i = 0; i < 30; i = i + 1) begin
            for (j = 0; j < 196; j = j + 1) begin
                weights_HL[(i * 196 + j) * 8 +: 8] = weights_HL_param[i * 196 + j];
            end
            biases_HL[i * 8 +: 8] = biases_HL_param[i];
        end
    end

endmodule
