/**********
* 1st dense layer implementation (output layer)
*
* Inputs: clk => clock signal, enable => enable signal, 
*         reset => active high sync reset, in_data => in vector, 
*
* Outputs: layer_out => dense layer output
*          layer_done => done signal
* 
***********/

module output_layer #(
  parameter HL_neurons = 32,
  parameter WIDTH = 8,
  parameter OL_neurons = 10
	)(
  input clk,
  input output_go,
  input reset,
  input signed [4*WIDTH*HL_neurons-1:0] output_in,
  output signed [4*WIDTH*OL_neurons-1:0] output_out,
  output output_done
  );
    
  wire signed [4*WIDTH*OL_neurons-1:0] dense_out;
  wire dense_done;

  //Biases and weights
  localparam signed [WIDTH*OL_neurons-1:0] biases_OL_param = { 8'sb11101111, 8'sb00001101, 8'sb11111100, 8'sb00000110, 8'sb00000011, 8'sb00000111, 8'sb11110111, 8'sb11111101, 8'sb11110110, 8'sb00001001 };
  
  localparam signed [WIDTH*HL_neurons*OL_neurons-1:0] weights_OL_param =  {
  8'sb11011000, 8'sb00001101, 8'sb11110111, 8'sb11111111, 8'sb11110000, 8'sb00001011, 8'sb00010000, 8'sb00010101, 8'sb11111100, 8'sb11111110, 8'sb11000100, 8'sb00010001, 8'sb00010111, 8'sb00010000, 8'sb11000000, 8'sb11100101, 8'sb00100011, 8'sb11011101, 8'sb00001011, 8'sb10111100, 8'sb11101101, 8'sb11000110, 8'sb11111100, 8'sb00010110, 8'sb00010011, 8'sb00000010, 8'sb11110111, 8'sb11101100, 8'sb00011111, 8'sb11111010, 8'sb00011001, 8'sb10111010,
  8'sb11111111, 8'sb10111110, 8'sb11001110, 8'sb11100111, 8'sb00001010, 8'sb11001110, 8'sb00010001, 8'sb00010111, 8'sb11101000, 8'sb11101010, 8'sb00001001, 8'sb00101010, 8'sb11010000, 8'sb00001110, 8'sb00101001, 8'sb10110001, 8'sb11011010, 8'sb11100011, 8'sb00010101, 8'sb00001111, 8'sb11110010, 8'sb00011110, 8'sb00011001, 8'sb11110100, 8'sb11110001, 8'sb00000001, 8'sb00011011, 8'sb10111100, 8'sb00100100, 8'sb00000001, 8'sb11011000, 8'sb00100101,
  8'sb01001001, 8'sb00000011, 8'sb11010111, 8'sb00100101, 8'sb00011011, 8'sb11100111, 8'sb11000111, 8'sb00000111, 8'sb00001011, 8'sb11111001, 8'sb11100001, 8'sb00101000, 8'sb00011100, 8'sb00000101, 8'sb00011111, 8'sb00100010, 8'sb00000011, 8'sb11101001, 8'sb11110101, 8'sb00011100, 8'sb11010011, 8'sb00000101, 8'sb11101001, 8'sb00001101, 8'sb10110100, 8'sb11101011, 8'sb11111010, 8'sb00011001, 8'sb00000010, 8'sb00000001, 8'sb00011010, 8'sb00001101,
  8'sb11110010, 8'sb11101000, 8'sb00000100, 8'sb11101110, 8'sb11111110, 8'sb11001110, 8'sb11011101, 8'sb11000011, 8'sb11111110, 8'sb11110010, 8'sb00100100, 8'sb00011010, 8'sb11110110, 8'sb11100101, 8'sb11001011, 8'sb00000010, 8'sb11100000, 8'sb11101101, 8'sb00000001, 8'sb11110100, 8'sb00001010, 8'sb00100011, 8'sb11101100, 8'sb11111011, 8'sb11100001, 8'sb00100101, 8'sb10100110, 8'sb00100110, 8'sb11110101, 8'sb00011010, 8'sb00011100, 8'sb11111000,
  8'sb10110110, 8'sb11111101, 8'sb00001011, 8'sb00110100, 8'sb11111110, 8'sb11111110, 8'sb00010000, 8'sb00010101, 8'sb11011110, 8'sb11001111, 8'sb00011101, 8'sb11011010, 8'sb10111011, 8'sb00110001, 8'sb00010001, 8'sb00001110, 8'sb10100111, 8'sb11111101, 8'sb11011001, 8'sb11110110, 8'sb00011100, 8'sb11101101, 8'sb11011100, 8'sb11110100, 8'sb00100010, 8'sb11001111, 8'sb00101111, 8'sb00001100, 8'sb11001011, 8'sb11101100, 8'sb00011011, 8'sb11011111,
  8'sb11110011, 8'sb11010000, 8'sb00011011, 8'sb00011010, 8'sb11100010, 8'sb11110010, 8'sb11111000, 8'sb10100101, 8'sb11010111, 8'sb01011100, 8'sb11111011, 8'sb10110111, 8'sb00011000, 8'sb11001001, 8'sb00000001, 8'sb11101011, 8'sb00010010, 8'sb00011000, 8'sb11101110, 8'sb00101010, 8'sb00010011, 8'sb00001000, 8'sb00011010, 8'sb00010111, 8'sb00010110, 8'sb00001101, 8'sb11101110, 8'sb00001101, 8'sb00001011, 8'sb11011111, 8'sb11110110, 8'sb00100011,
  8'sb11101101, 8'sb00010000, 8'sb11111111, 8'sb11101000, 8'sb00001001, 8'sb00110010, 8'sb00100110, 8'sb11111001, 8'sb10111001, 8'sb11001110, 8'sb10110110, 8'sb10111110, 8'sb00010001, 8'sb11110000, 8'sb00010111, 8'sb00011100, 8'sb00101111, 8'sb10110111, 8'sb11101110, 8'sb00001100, 8'sb11101000, 8'sb00010000, 8'sb00011101, 8'sb00011001, 8'sb00001011, 8'sb11101011, 8'sb00011001, 8'sb11001010, 8'sb11101000, 8'sb11100111, 8'sb11111010, 8'sb11101001,
  8'sb00001111, 8'sb11110010, 8'sb00000111, 8'sb10111011, 8'sb11111010, 8'sb11010101, 8'sb11100100, 8'sb00011101, 8'sb00001101, 8'sb00001000, 8'sb11111101, 8'sb00101111, 8'sb10111111, 8'sb00010100, 8'sb11001101, 8'sb00000001, 8'sb11110011, 8'sb00010011, 8'sb11001111, 8'sb11110011, 8'sb11110001, 8'sb11011011, 8'sb00100111, 8'sb10101101, 8'sb00101100, 8'sb11101001, 8'sb00001110, 8'sb00100101, 8'sb00100100, 8'sb00000110, 8'sb00001001, 8'sb00111001,
  8'sb11100100, 8'sb00000001, 8'sb00000111, 8'sb00011010, 8'sb00000011, 8'sb00010111, 8'sb11000010, 8'sb00000111, 8'sb00010000, 8'sb11101110, 8'sb00000010, 8'sb11011100, 8'sb00001111, 8'sb00001001, 8'sb11111101, 8'sb11110001, 8'sb00010010, 8'sb00011110, 8'sb00010010, 8'sb11111000, 8'sb11110101, 8'sb00001111, 8'sb11011000, 8'sb00001000, 8'sb11101110, 8'sb00000010, 8'sb00011110, 8'sb11011001, 8'sb10110110, 8'sb00010011, 8'sb11011001, 8'sb11011110,
  8'sb10000001, 8'sb00010000, 8'sb00000101, 8'sb10110011, 8'sb10011011, 8'sb11111000, 8'sb00001100, 8'sb00001100, 8'sb00011001, 8'sb00001011, 8'sb00010000, 8'sb11110101, 8'sb00000000, 8'sb11010101, 8'sb00010101, 8'sb00010101, 8'sb11101000, 8'sb11110100, 8'sb00010011, 8'sb00001010, 8'sb00011100, 8'sb11101011, 8'sb11010100, 8'sb11011111, 8'sb00011001, 8'sb11110000, 8'sb10111110, 8'sb00010010, 8'sb11111111, 8'sb00100011, 8'sb11000100, 8'sb10011011
  };
  
  dense_layer #(
    .NEURON_NB(OL_neurons),
    .IN_SIZE(HL_neurons), 
    .WIDTH(WIDTH),
    .WIDTH_IN(4*WIDTH),
    .WIDTH_OUT(4*WIDTH)
  ) output_dense (
    .clk(clk), 
    .dense_go(output_go), 
    .reset(reset),
    .dense_in(output_in), 
    .weights(weights_OL_param), 
    .biases(biases_OL_param),
    .dense_out(dense_out), 
    .dense_done(dense_done)
  ); //Dense layer

  ReLU_layer #(
    .NEURON_NB(OL_neurons),
    .IN_SIZE(HL_neurons),
    .WIDTH(4*WIDTH)
  ) ReLU_output_layer (
    .clk(clk),
    .reset(reset),
    .relu_go(dense_done),
    .data_in_array(dense_out),
    .relu_layer_done(output_done),
    .data_out_array(output_out)
  );

endmodule
