module MLP #(
    //constants
    parameter averaged_pixels_nr = 196,
    parameter resolution = 8,
    parameter HL_neurons = 30,
    parameter OL_neurons = 10
	)(
    input clk,
    input reset,
    input signed [resolution*averaged_pixels_nr-1:0] averaged_pixels,
    output signed [resolution*OL_neurons-1:0] output_activations
    );

    // Intermediate signals
    wire signed [resolution*HL_neurons-1:0] zeds_HL;
    wire signed [resolution*HL_neurons-1:0] activations_HL;
    wire signed [resolution*HL_neurons-1:0] activations_HL_w;
    wire signed [resolution*OL_neurons-1:0] zeds_OL;
    wire signed [resolution*OL_neurons-1:0] activations_OL;

    // Local parameters for initialized weights and biases
    localparam signed [8*30*196-1:0] weights_HL_param = {
    8'sb00001011, 8'sb00001010, 8'sb00001011, 8'sb00001011, 8'sb00001100, 8'sb00001011, 8'sb00001110, 8'sb00001101, 8'sb00001011, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00001110, 8'sb00001100, 8'sb00001010, 8'sb00001010, 8'sb00001011, 8'sb00001101, 8'sb00010000, 8'sb00010001, 8'sb00010101, 8'sb00010010, 8'sb00010001, 8'sb00010001, 8'sb00010000, 8'sb00010001, 8'sb00001101, 8'sb00001010, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00001101, 8'sb00001001, 8'sb00010010, 8'sb00010111, 8'sb00011001, 8'sb00010111, 8'sb00011001, 8'sb00010100, 8'sb00001011, 8'sb00001101, 8'sb00001111, 8'sb00001110, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00001101, 8'sb00010000, 8'sb00010001, 8'sb00010101, 8'sb00001000, 8'sb00011000, 8'sb00010011, 8'sb00010000, 8'sb00010110, 8'sb00001101, 8'sb00001101, 8'sb00001100, 8'sb00001110, 8'sb00001111, 8'sb00001111, 8'sb00001011, 8'sb00001001, 8'sb00001101, 8'sb00010110, 8'sb00001111, 8'sb00011000, 8'sb00011010, 8'sb00100011, 8'sb00010010, 8'sb00001100, 8'sb00001110, 8'sb00001111, 8'sb00001000, 8'sb00000110, 8'sb00001101, 8'sb00001000, 8'sb00010011, 8'sb11111000, 8'sb11111111, 8'sb00001011, 8'sb00100000, 8'sb00100100, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00001010, 8'sb00001010, 8'sb00000010, 8'sb00011100, 8'sb00000100, 8'sb11110110, 8'sb11111111, 8'sb00000011, 8'sb00010111, 8'sb00010011, 8'sb00001011, 8'sb00001011, 8'sb00001110, 8'sb00000100, 8'sb00000011, 8'sb00001000, 8'sb00010000, 8'sb00011011, 8'sb00001010, 8'sb11111000, 8'sb11110001, 8'sb00000111, 8'sb00001010, 8'sb00001110, 8'sb00001001, 8'sb00001101, 8'sb00001110, 8'sb00000000, 8'sb11111100, 8'sb00001010, 8'sb00010100, 8'sb00011010, 8'sb11111010, 8'sb11110110, 8'sb11111100, 8'sb00001000, 8'sb00010011, 8'sb00001100, 8'sb00001010, 8'sb00001100, 8'sb00001101, 8'sb00001100, 8'sb00011100, 8'sb00010110, 8'sb00010010, 8'sb00001111, 8'sb11111100, 8'sb00010001, 8'sb00011010, 8'sb00010110, 8'sb00010101, 8'sb00001010, 8'sb00001010, 8'sb00001110, 8'sb00010000, 8'sb00011001, 8'sb00100111, 8'sb00100100, 8'sb00101010, 8'sb00110011, 8'sb00110010, 8'sb00101000, 8'sb00101111, 8'sb00101000, 8'sb00010101, 8'sb00000111, 8'sb00001011, 8'sb00001110, 8'sb00001110, 8'sb00010111, 8'sb00010100, 8'sb00011000, 8'sb00010111, 8'sb00100100, 8'sb00011110, 8'sb00100100, 8'sb00100110, 8'sb00100001, 8'sb00001101, 8'sb00001011, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00000110, 8'sb00001000, 8'sb00010101, 8'sb00010110, 8'sb00011101, 8'sb00011111, 8'sb00011100, 8'sb00010100, 8'sb00000111, 8'sb00001010, 8'sb00001100, 8'sb00001011, 8'sb00001010, 8'sb00001010, 8'sb00001100, 8'sb00001100, 8'sb00000111, 8'sb00001010, 8'sb00001011, 8'sb00001000, 8'sb00001100, 8'sb00001001, 8'sb00001100, 8'sb00001110, 8'sb00001101, 8'sb00001010,
    8'sb00001011, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001011, 8'sb00001100, 8'sb00001010, 8'sb00001011, 8'sb00001110, 8'sb00001010, 8'sb00001100, 8'sb00001101, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00001101, 8'sb00001010, 8'sb00001100, 8'sb00001001, 8'sb00001010, 8'sb00010010, 8'sb00001110, 8'sb00000110, 8'sb00000011, 8'sb00000111, 8'sb00000100, 8'sb00001010, 8'sb00001101, 8'sb00001100, 8'sb00001101, 8'sb00001100, 8'sb00010000, 8'sb00010100, 8'sb00011010, 8'sb00011001, 8'sb00011010, 8'sb00100100, 8'sb00011111, 8'sb00001010, 8'sb00000001, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001100, 8'sb00010100, 8'sb00011000, 8'sb00001111, 8'sb00010001, 8'sb00010101, 8'sb00001100, 8'sb00001011, 8'sb00011111, 8'sb00011011, 8'sb00011000, 8'sb00010110, 8'sb00001101, 8'sb00001101, 8'sb00001010, 8'sb00010010, 8'sb00010010, 8'sb00010010, 8'sb00100010, 8'sb00100000, 8'sb00010011, 8'sb00010010, 8'sb00011010, 8'sb00011001, 8'sb00100010, 8'sb00100011, 8'sb00010010, 8'sb00001101, 8'sb00001100, 8'sb00001110, 8'sb00001011, 8'sb00000100, 8'sb00000111, 8'sb00010001, 8'sb00010001, 8'sb00000000, 8'sb00001110, 8'sb00001110, 8'sb00010011, 8'sb00100000, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00000110, 8'sb00000101, 8'sb00000100, 8'sb11111110, 8'sb00011110, 8'sb00010000, 8'sb00000011, 8'sb00001101, 8'sb11111100, 8'sb11110100, 8'sb00000010, 8'sb00001101, 8'sb00001010, 8'sb00001100, 8'sb00001011, 8'sb00000111, 8'sb00001110, 8'sb00000011, 8'sb00010101, 8'sb00001000, 8'sb11111100, 8'sb11111101, 8'sb11111010, 8'sb00000010, 8'sb00001001, 8'sb00010000, 8'sb00001100, 8'sb00010000, 8'sb00010101, 8'sb11111110, 8'sb00000100, 8'sb00001010, 8'sb00001110, 8'sb00000000, 8'sb00000101, 8'sb00001010, 8'sb00010011, 8'sb00011011, 8'sb00010100, 8'sb00001100, 8'sb00001100, 8'sb00001111, 8'sb00011110, 8'sb00010001, 8'sb00010000, 8'sb00010001, 8'sb00000000, 8'sb00011001, 8'sb00011011, 8'sb00011010, 8'sb00011010, 8'sb00100111, 8'sb00010111, 8'sb00001110, 8'sb00001011, 8'sb00001111, 8'sb00011011, 8'sb00100101, 8'sb00010011, 8'sb00010000, 8'sb00000101, 8'sb00010000, 8'sb00010011, 8'sb00010001, 8'sb00100001, 8'sb00100001, 8'sb00010000, 8'sb00001100, 8'sb00001010, 8'sb00010000, 8'sb00010100, 8'sb00011101, 8'sb00001101, 8'sb00010000, 8'sb00001110, 8'sb00000111, 8'sb00010101, 8'sb00010001, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00001101, 8'sb00001010, 8'sb00001110, 8'sb00001001, 8'sb00000101, 8'sb00010010, 8'sb00010100, 8'sb00011000, 8'sb00010101, 8'sb00010110, 8'sb00001110, 8'sb00000101, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00001011, 8'sb00001100, 8'sb00001100, 8'sb00001101, 8'sb00010000, 8'sb00010010, 8'sb00010011, 8'sb00001011, 8'sb00001001, 8'sb00001100, 8'sb00001100, 8'sb00001101,
    8'sb00010001, 8'sb00001101, 8'sb00001111, 8'sb00010001, 8'sb00001101, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00001111, 8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00001100, 8'sb00001100, 8'sb00010001, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010011, 8'sb00010101, 8'sb00011010, 8'sb00010101, 8'sb00010111, 8'sb00010011, 8'sb00001110, 8'sb00001100, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00010001, 8'sb00010100, 8'sb00011101, 8'sb00100100, 8'sb00011010, 8'sb00010011, 8'sb00010011, 8'sb00010100, 8'sb00010101, 8'sb00001010, 8'sb00001010, 8'sb00001101, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00011100, 8'sb00100100, 8'sb00010111, 8'sb00001111, 8'sb00010111, 8'sb00001011, 8'sb00001110, 8'sb00001111, 8'sb00001001, 8'sb00000100, 8'sb00000010, 8'sb00001101, 8'sb00010000, 8'sb00010010, 8'sb00100000, 8'sb00001000, 8'sb00000000, 8'sb00000000, 8'sb00001000, 8'sb00010111, 8'sb00100001, 8'sb00001110, 8'sb00001101, 8'sb00000100, 8'sb11110111, 8'sb00001001, 8'sb00001100, 8'sb00010010, 8'sb00000110, 8'sb11100010, 8'sb11101101, 8'sb11110001, 8'sb11111011, 8'sb11110110, 8'sb00011011, 8'sb00010011, 8'sb00010110, 8'sb00010000, 8'sb00000011, 8'sb00001011, 8'sb00010000, 8'sb00001110, 8'sb11111111, 8'sb00000100, 8'sb00001111, 8'sb00001100, 8'sb00001111, 8'sb11110110, 8'sb00010010, 8'sb11111110, 8'sb00000000, 8'sb00100100, 8'sb00100010, 8'sb00001110, 8'sb00001110, 8'sb00001111, 8'sb00011001, 8'sb00100000, 8'sb00011001, 8'sb00010001, 8'sb00000111, 8'sb11110101, 8'sb00010000, 8'sb00001010, 8'sb00011000, 8'sb00100011, 8'sb00011010, 8'sb00001111, 8'sb00001100, 8'sb00010001, 8'sb00010001, 8'sb00011100, 8'sb00011101, 8'sb00010000, 8'sb00001001, 8'sb00001000, 8'sb00011110, 8'sb00011111, 8'sb00011110, 8'sb00100000, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00010110, 8'sb00001101, 8'sb00010000, 8'sb00010000, 8'sb00010010, 8'sb00001000, 8'sb00010111, 8'sb00011110, 8'sb00011010, 8'sb00011001, 8'sb00010010, 8'sb00001100, 8'sb00010001, 8'sb00010000, 8'sb00010101, 8'sb00010011, 8'sb00010111, 8'sb00010001, 8'sb00010110, 8'sb00010111, 8'sb00010010, 8'sb00010100, 8'sb00010110, 8'sb00010101, 8'sb00000011, 8'sb00001101, 8'sb00001111, 8'sb00001101, 8'sb00010011, 8'sb00010000, 8'sb00010010, 8'sb00010000, 8'sb00010101, 8'sb00001111, 8'sb00010001, 8'sb00000111, 8'sb00001010, 8'sb00000101, 8'sb00001001, 8'sb00001101, 8'sb00001100, 8'sb00001110, 8'sb00010000, 8'sb00010110, 8'sb00011001, 8'sb00011001, 8'sb00010110, 8'sb00010011, 8'sb00001110, 8'sb00001111, 8'sb00000000, 8'sb00000010, 8'sb00001011, 8'sb00010000, 8'sb00010001, 8'sb00001100, 8'sb00010001, 8'sb00001101, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00010000, 8'sb00001101, 8'sb00010000, 8'sb00001111, 8'sb00001110, 8'sb00001111, 8'sb00001110,
    8'sb00001111, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00010011, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010011, 8'sb00001111, 8'sb00001111, 8'sb00010000, 8'sb00001101, 8'sb00001110, 8'sb00001111, 8'sb00010001, 8'sb00010010, 8'sb00001111, 8'sb00010010, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00010100, 8'sb00010001, 8'sb00001101, 8'sb00010110, 8'sb00010000, 8'sb00001101, 8'sb00001111, 8'sb00001101, 8'sb00010000, 8'sb00011000, 8'sb00010110, 8'sb00010010, 8'sb00010010, 8'sb00010010, 8'sb00010111, 8'sb00001101, 8'sb00010100, 8'sb00010010, 8'sb00010100, 8'sb00010010, 8'sb00010101, 8'sb00010010, 8'sb00010100, 8'sb00010010, 8'sb00011110, 8'sb00010101, 8'sb00010010, 8'sb00010101, 8'sb00010100, 8'sb00010000, 8'sb00011001, 8'sb00010011, 8'sb00010011, 8'sb00001110, 8'sb00001101, 8'sb00001010, 8'sb00001011, 8'sb00001101, 8'sb00011101, 8'sb00010100, 8'sb00010011, 8'sb00010110, 8'sb00001101, 8'sb00000111, 8'sb00000110, 8'sb00000100, 8'sb00001101, 8'sb11111111, 8'sb00000010, 8'sb00000110, 8'sb00000000, 8'sb11111011, 8'sb00001011, 8'sb00010001, 8'sb00010011, 8'sb00010110, 8'sb00010001, 8'sb00001001, 8'sb00010000, 8'sb00001111, 8'sb00010110, 8'sb00001110, 8'sb00010000, 8'sb00001100, 8'sb00000100, 8'sb11111100, 8'sb00000011, 8'sb00001111, 8'sb00010000, 8'sb00010000, 8'sb00001101, 8'sb00000110, 8'sb00011000, 8'sb00010110, 8'sb00010111, 8'sb00010001, 8'sb00000101, 8'sb00001001, 8'sb00010000, 8'sb00011000, 8'sb00001110, 8'sb00010000, 8'sb00010011, 8'sb00010100, 8'sb11111010, 8'sb11011011, 8'sb11101000, 8'sb00001010, 8'sb00011100, 8'sb00000100, 8'sb00001010, 8'sb00011000, 8'sb00010010, 8'sb00011010, 8'sb00010100, 8'sb00010001, 8'sb00010010, 8'sb00011001, 8'sb00000001, 8'sb11101110, 8'sb11011100, 8'sb11000010, 8'sb11001001, 8'sb11111011, 8'sb00001110, 8'sb00010001, 8'sb00010001, 8'sb00010011, 8'sb00010001, 8'sb00010001, 8'sb00010010, 8'sb00010111, 8'sb00010110, 8'sb00001110, 8'sb00010111, 8'sb00100001, 8'sb00100000, 8'sb00010100, 8'sb00001000, 8'sb00001011, 8'sb00010000, 8'sb00001100, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00010010, 8'sb00011100, 8'sb00011011, 8'sb00010111, 8'sb00011110, 8'sb00011100, 8'sb00011100, 8'sb00010011, 8'sb00010010, 8'sb00001001, 8'sb00001111, 8'sb00001111, 8'sb00010010, 8'sb00010000, 8'sb00010001, 8'sb00011000, 8'sb00101001, 8'sb00100101, 8'sb00011110, 8'sb00011000, 8'sb00010011, 8'sb00010001, 8'sb00001011, 8'sb00010000, 8'sb00010101, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00010001, 8'sb00010000, 8'sb00010100, 8'sb00010001, 8'sb00010110, 8'sb00010100, 8'sb00010010, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00010011,
    8'sb00001010, 8'sb00001100, 8'sb00001011, 8'sb00001011, 8'sb00001011, 8'sb00001100, 8'sb00001100, 8'sb00001101, 8'sb00001110, 8'sb00001011, 8'sb00001011, 8'sb00001100, 8'sb00001111, 8'sb00001100, 8'sb00001010, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00001011, 8'sb00001011, 8'sb00001011, 8'sb00001101, 8'sb00001101, 8'sb00010001, 8'sb00010001, 8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00001011, 8'sb00001011, 8'sb00001111, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00001001, 8'sb00000100, 8'sb00001000, 8'sb00010011, 8'sb00010001, 8'sb00010001, 8'sb00010000, 8'sb00001101, 8'sb00001100, 8'sb00001011, 8'sb00010011, 8'sb00010011, 8'sb00010101, 8'sb00010011, 8'sb00010000, 8'sb00001101, 8'sb00001111, 8'sb00011101, 8'sb00001111, 8'sb00001110, 8'sb00010010, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00010000, 8'sb00010010, 8'sb00001011, 8'sb00001110, 8'sb00001001, 8'sb00001011, 8'sb00001100, 8'sb00001110, 8'sb00011100, 8'sb00011001, 8'sb00011001, 8'sb00001111, 8'sb00001010, 8'sb00001100, 8'sb00010000, 8'sb00010001, 8'sb00001001, 8'sb00001101, 8'sb00001110, 8'sb00001101, 8'sb00100000, 8'sb00000100, 8'sb11111101, 8'sb00000010, 8'sb00001000, 8'sb00001110, 8'sb00001100, 8'sb00001111, 8'sb00011011, 8'sb00010111, 8'sb00010011, 8'sb00010110, 8'sb00001101, 8'sb00010100, 8'sb00100101, 8'sb00011100, 8'sb00001010, 8'sb11111000, 8'sb11111110, 8'sb00001010, 8'sb00001110, 8'sb00001110, 8'sb00001111, 8'sb00000100, 8'sb11111001, 8'sb11111110, 8'sb00000100, 8'sb00011011, 8'sb00011011, 8'sb00011000, 8'sb00011101, 8'sb00010000, 8'sb00000101, 8'sb00001011, 8'sb00001100, 8'sb00001111, 8'sb00000101, 8'sb00000101, 8'sb00000000, 8'sb11100110, 8'sb00001111, 8'sb00100001, 8'sb00001110, 8'sb00011001, 8'sb00010100, 8'sb00000110, 8'sb00000100, 8'sb00001011, 8'sb00001100, 8'sb00010011, 8'sb00001111, 8'sb00001111, 8'sb00000010, 8'sb11101011, 8'sb00100001, 8'sb00011101, 8'sb00011000, 8'sb00010111, 8'sb00010000, 8'sb11111110, 8'sb00000001, 8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00001101, 8'sb00000010, 8'sb11111101, 8'sb11111100, 8'sb00001111, 8'sb00011010, 8'sb00101001, 8'sb00010110, 8'sb00001111, 8'sb00001001, 8'sb00001010, 8'sb00001011, 8'sb00001100, 8'sb00001011, 8'sb00001111, 8'sb11111100, 8'sb11111110, 8'sb00000110, 8'sb11111101, 8'sb00001111, 8'sb00010111, 8'sb00010110, 8'sb00010010, 8'sb00010001, 8'sb00001111, 8'sb00001101, 8'sb00001011, 8'sb00001110, 8'sb00010111, 8'sb00100010, 8'sb00011000, 8'sb00001100, 8'sb00001010, 8'sb00010010, 8'sb00010110, 8'sb00010111, 8'sb00010111, 8'sb00010011, 8'sb00001010, 8'sb00001100, 8'sb00001011, 8'sb00001110, 8'sb00001101, 8'sb00010000, 8'sb00010010, 8'sb00010000, 8'sb00010010, 8'sb00010001, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001100, 8'sb00001101,
    8'sb00010100, 8'sb00010011, 8'sb00010011, 8'sb00010011, 8'sb00010000, 8'sb00010001, 8'sb00010000, 8'sb00010100, 8'sb00010000, 8'sb00010000, 8'sb00010011, 8'sb00010100, 8'sb00010000, 8'sb00010100, 8'sb00010010, 8'sb00010011, 8'sb00010001, 8'sb00010011, 8'sb00010111, 8'sb00011010, 8'sb00011000, 8'sb00010001, 8'sb00010000, 8'sb00001101, 8'sb00001011, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00010100, 8'sb00010011, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00011000, 8'sb00001100, 8'sb00001010, 8'sb00001000, 8'sb00010000, 8'sb00010100, 8'sb00010100, 8'sb00010010, 8'sb00001101, 8'sb00000001, 8'sb00000110, 8'sb00001110, 8'sb00000111, 8'sb00010100, 8'sb00010100, 8'sb00010000, 8'sb00010001, 8'sb00001010, 8'sb00000100, 8'sb00010010, 8'sb00010001, 8'sb00010000, 8'sb00001101, 8'sb00001010, 8'sb00010001, 8'sb00011001, 8'sb00000110, 8'sb00001001, 8'sb00010000, 8'sb00001001, 8'sb00001000, 8'sb11111101, 8'sb11111101, 8'sb00010100, 8'sb00010001, 8'sb00010000, 8'sb00001001, 8'sb11111110, 8'sb00000110, 8'sb11111110, 8'sb11110100, 8'sb00000110, 8'sb00011010, 8'sb00000110, 8'sb00001100, 8'sb11111100, 8'sb00001101, 8'sb00010010, 8'sb00010011, 8'sb00010010, 8'sb11110111, 8'sb11011111, 8'sb11100101, 8'sb11110011, 8'sb00000001, 8'sb00000001, 8'sb00000111, 8'sb00000111, 8'sb00010000, 8'sb00000000, 8'sb00001110, 8'sb00010101, 8'sb00010010, 8'sb00010100, 8'sb00000101, 8'sb00001101, 8'sb00011100, 8'sb00011110, 8'sb00011101, 8'sb00001010, 8'sb00000101, 8'sb11110110, 8'sb11110110, 8'sb00000100, 8'sb00011000, 8'sb00011000, 8'sb00010001, 8'sb00010011, 8'sb00011100, 8'sb00011101, 8'sb00010111, 8'sb00010110, 8'sb00101010, 8'sb00010000, 8'sb11111110, 8'sb00000000, 8'sb00010010, 8'sb00011011, 8'sb00100110, 8'sb00010111, 8'sb00010010, 8'sb00001111, 8'sb00011001, 8'sb00010110, 8'sb00011101, 8'sb00011101, 8'sb00101001, 8'sb11110001, 8'sb00000001, 8'sb00001100, 8'sb00010110, 8'sb00011001, 8'sb00100111, 8'sb00010110, 8'sb00010001, 8'sb00010010, 8'sb00011011, 8'sb00010000, 8'sb00010110, 8'sb00011000, 8'sb00000111, 8'sb00000000, 8'sb00001010, 8'sb00010110, 8'sb00001000, 8'sb00010111, 8'sb00011100, 8'sb00010011, 8'sb00010010, 8'sb00010001, 8'sb00011010, 8'sb00001110, 8'sb00001100, 8'sb00001000, 8'sb00001111, 8'sb00000110, 8'sb00001010, 8'sb00011010, 8'sb00010110, 8'sb00010101, 8'sb00010011, 8'sb00010011, 8'sb00010100, 8'sb00010001, 8'sb00001101, 8'sb00000010, 8'sb11111110, 8'sb00000011, 8'sb00001110, 8'sb00001101, 8'sb00001011, 8'sb00001001, 8'sb00010000, 8'sb00010001, 8'sb00010100, 8'sb00010101, 8'sb00010100, 8'sb00010011, 8'sb00010101, 8'sb00001111, 8'sb00010001, 8'sb00010001, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00010100, 8'sb00010001, 8'sb00010010,
    8'sb00010100, 8'sb00010010, 8'sb00010011, 8'sb00010000, 8'sb00010100, 8'sb00010000, 8'sb00010010, 8'sb00010000, 8'sb00010000, 8'sb00010100, 8'sb00010001, 8'sb00010010, 8'sb00010011, 8'sb00010101, 8'sb00010100, 8'sb00010100, 8'sb00010010, 8'sb00010000, 8'sb00001111, 8'sb00001010, 8'sb00000111, 8'sb00000010, 8'sb00000101, 8'sb00001101, 8'sb00001100, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00010101, 8'sb00010001, 8'sb00000111, 8'sb11111110, 8'sb11111011, 8'sb11111101, 8'sb00000000, 8'sb11111001, 8'sb11111010, 8'sb00000001, 8'sb00001010, 8'sb00001110, 8'sb00010011, 8'sb00010101, 8'sb00010011, 8'sb00010101, 8'sb00001011, 8'sb00001001, 8'sb00001000, 8'sb00000011, 8'sb00001110, 8'sb00010001, 8'sb00001110, 8'sb00010101, 8'sb00011010, 8'sb00011100, 8'sb00010011, 8'sb00010010, 8'sb00011001, 8'sb00010110, 8'sb00010001, 8'sb00010001, 8'sb11111011, 8'sb00010101, 8'sb00010101, 8'sb00100001, 8'sb00011100, 8'sb00010111, 8'sb00011010, 8'sb00100000, 8'sb00010110, 8'sb00010001, 8'sb00010111, 8'sb00001100, 8'sb00000001, 8'sb00001110, 8'sb00100000, 8'sb00010010, 8'sb00010100, 8'sb00010110, 8'sb00001101, 8'sb00010001, 8'sb00011110, 8'sb00100011, 8'sb00010110, 8'sb00010101, 8'sb00010110, 8'sb00010010, 8'sb00011111, 8'sb00100001, 8'sb00011001, 8'sb00000001, 8'sb00010010, 8'sb00010000, 8'sb00000010, 8'sb11111110, 8'sb11111100, 8'sb00001011, 8'sb00010011, 8'sb00010010, 8'sb00010110, 8'sb00010000, 8'sb00010001, 8'sb00010110, 8'sb00000110, 8'sb00001000, 8'sb00010000, 8'sb00100101, 8'sb00001110, 8'sb00001110, 8'sb00000111, 8'sb00001010, 8'sb00010011, 8'sb00010001, 8'sb00001101, 8'sb11111111, 8'sb00000101, 8'sb00010100, 8'sb00010010, 8'sb00010111, 8'sb00010101, 8'sb00001011, 8'sb00000110, 8'sb00001100, 8'sb11111100, 8'sb00000001, 8'sb00001111, 8'sb00010011, 8'sb00001110, 8'sb11110010, 8'sb11111011, 8'sb00000110, 8'sb00001101, 8'sb00011011, 8'sb00001110, 8'sb11111011, 8'sb00000101, 8'sb00000001, 8'sb11110000, 8'sb00000010, 8'sb00010011, 8'sb00010010, 8'sb00001110, 8'sb11110100, 8'sb11111100, 8'sb00000010, 8'sb11111100, 8'sb00000100, 8'sb00001011, 8'sb00000010, 8'sb11111110, 8'sb11111111, 8'sb00000101, 8'sb00001100, 8'sb00010001, 8'sb00010001, 8'sb00001111, 8'sb00001101, 8'sb00001110, 8'sb00001111, 8'sb00010000, 8'sb00001010, 8'sb00001100, 8'sb00001000, 8'sb00000100, 8'sb00000001, 8'sb00010001, 8'sb00010010, 8'sb00010100, 8'sb00010100, 8'sb00010101, 8'sb00010001, 8'sb00010101, 8'sb00010001, 8'sb00001101, 8'sb00001010, 8'sb00010001, 8'sb00001010, 8'sb00010010, 8'sb00010001, 8'sb00010101, 8'sb00010000, 8'sb00010100, 8'sb00010001, 8'sb00010001, 8'sb00010101, 8'sb00010100, 8'sb00010011, 8'sb00010100, 8'sb00010100, 8'sb00010111, 8'sb00010001, 8'sb00010011, 8'sb00010001, 8'sb00010100, 8'sb00010001, 8'sb00010010,
    8'sb00001111, 8'sb00010001, 8'sb00010001, 8'sb00010011, 8'sb00010001, 8'sb00010100, 8'sb00010100, 8'sb00010011, 8'sb00010001, 8'sb00010000, 8'sb00010000, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00010001, 8'sb00010001, 8'sb00010010, 8'sb00010001, 8'sb00011000, 8'sb00010110, 8'sb00010101, 8'sb00011010, 8'sb00010011, 8'sb00010001, 8'sb00001101, 8'sb00010000, 8'sb00010001, 8'sb00010011, 8'sb00010011, 8'sb00010011, 8'sb00010000, 8'sb00010010, 8'sb00001111, 8'sb00001110, 8'sb00011000, 8'sb00011000, 8'sb00000101, 8'sb00000011, 8'sb00001010, 8'sb00001101, 8'sb00001111, 8'sb00010001, 8'sb00010010, 8'sb00010011, 8'sb00010000, 8'sb00011001, 8'sb00001101, 8'sb00001110, 8'sb00000101, 8'sb11110100, 8'sb00001001, 8'sb00001010, 8'sb00000111, 8'sb00000100, 8'sb00001010, 8'sb00001110, 8'sb00010100, 8'sb00011010, 8'sb00011001, 8'sb00010111, 8'sb00001111, 8'sb00010010, 8'sb00001011, 8'sb00001010, 8'sb00001000, 8'sb00001100, 8'sb00001011, 8'sb00001110, 8'sb00000111, 8'sb00001111, 8'sb00010010, 8'sb00011100, 8'sb00011011, 8'sb00010010, 8'sb00010010, 8'sb00011011, 8'sb00001101, 8'sb00001000, 8'sb00001101, 8'sb00001101, 8'sb00010010, 8'sb00010000, 8'sb00001101, 8'sb00001110, 8'sb00010010, 8'sb00011011, 8'sb00011010, 8'sb00011001, 8'sb00011101, 8'sb00001011, 8'sb11100011, 8'sb00001010, 8'sb00000110, 8'sb00010000, 8'sb00001100, 8'sb00010011, 8'sb00010101, 8'sb00010000, 8'sb00010000, 8'sb00010011, 8'sb00001011, 8'sb00001110, 8'sb00000101, 8'sb11011111, 8'sb00000001, 8'sb00010101, 8'sb00000110, 8'sb00001101, 8'sb00001110, 8'sb00011101, 8'sb00010110, 8'sb00010000, 8'sb00001111, 8'sb00001110, 8'sb00000110, 8'sb00000010, 8'sb11100101, 8'sb11011101, 8'sb00100010, 8'sb00011110, 8'sb00010101, 8'sb00001110, 8'sb00010010, 8'sb00001110, 8'sb00011000, 8'sb00010000, 8'sb00010011, 8'sb00010000, 8'sb00000100, 8'sb11110101, 8'sb11101010, 8'sb11111101, 8'sb00111011, 8'sb00011110, 8'sb00010100, 8'sb00010100, 8'sb00000110, 8'sb00001000, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00010000, 8'sb00000010, 8'sb11111101, 8'sb11111100, 8'sb00010110, 8'sb00100100, 8'sb00100100, 8'sb00010111, 8'sb00010101, 8'sb00000010, 8'sb00001010, 8'sb00010010, 8'sb00010100, 8'sb00010000, 8'sb00010001, 8'sb00001101, 8'sb00001010, 8'sb00000110, 8'sb11111100, 8'sb00001000, 8'sb00010000, 8'sb00011011, 8'sb00011001, 8'sb00001000, 8'sb00001001, 8'sb00010010, 8'sb00010010, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00001011, 8'sb00001010, 8'sb00000101, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00001100, 8'sb00001101, 8'sb00010001, 8'sb00001111, 8'sb00010011, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00010100, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00010010, 8'sb00011001, 8'sb00010100, 8'sb00010011, 8'sb00010001, 8'sb00010001,
    8'sb00001111, 8'sb00001101, 8'sb00001101, 8'sb00001011, 8'sb00001011, 8'sb00001100, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00001011, 8'sb00010000, 8'sb00001100, 8'sb00001110, 8'sb00001111, 8'sb00001110, 8'sb00000111, 8'sb11111111, 8'sb00000010, 8'sb11111110, 8'sb00001001, 8'sb00010100, 8'sb00001111, 8'sb00001011, 8'sb00001011, 8'sb00001100, 8'sb00001110, 8'sb00010000, 8'sb00010000, 8'sb00010001, 8'sb00001011, 8'sb00001100, 8'sb00001101, 8'sb00010011, 8'sb00000011, 8'sb11111111, 8'sb00000001, 8'sb00010010, 8'sb00011001, 8'sb00010101, 8'sb00010001, 8'sb00001100, 8'sb00001101, 8'sb00010110, 8'sb00010100, 8'sb00011000, 8'sb00011001, 8'sb00010111, 8'sb00011011, 8'sb00011101, 8'sb00011100, 8'sb00011101, 8'sb00101001, 8'sb00010101, 8'sb00001101, 8'sb00001111, 8'sb00010010, 8'sb00010000, 8'sb00010001, 8'sb00010100, 8'sb00010000, 8'sb00011101, 8'sb00011111, 8'sb00110000, 8'sb00100101, 8'sb00011010, 8'sb00011100, 8'sb00001101, 8'sb00001010, 8'sb00001111, 8'sb00010001, 8'sb00001110, 8'sb00010011, 8'sb00010111, 8'sb00011001, 8'sb00010101, 8'sb00001000, 8'sb00001111, 8'sb00001100, 8'sb00011000, 8'sb00010010, 8'sb00001101, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00011001, 8'sb00101011, 8'sb00100111, 8'sb00100010, 8'sb00010100, 8'sb00000011, 8'sb00001011, 8'sb00010010, 8'sb00001110, 8'sb00010110, 8'sb00001110, 8'sb00001111, 8'sb00001111, 8'sb00001100, 8'sb00011110, 8'sb00010110, 8'sb00011000, 8'sb00010100, 8'sb00000101, 8'sb00000111, 8'sb00010000, 8'sb00010010, 8'sb00001000, 8'sb00001110, 8'sb00001000, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00000011, 8'sb00001000, 8'sb00010111, 8'sb00010000, 8'sb00010010, 8'sb00000101, 8'sb00010110, 8'sb00010001, 8'sb00001110, 8'sb00010010, 8'sb00000010, 8'sb00001101, 8'sb00010000, 8'sb00001011, 8'sb11111110, 8'sb00000110, 8'sb11111111, 8'sb00000000, 8'sb11111111, 8'sb11111101, 8'sb00001010, 8'sb00001101, 8'sb00001000, 8'sb00001000, 8'sb11111110, 8'sb00001111, 8'sb00001111, 8'sb00001101, 8'sb00000000, 8'sb11111101, 8'sb11111000, 8'sb11110111, 8'sb11111101, 8'sb11111111, 8'sb00000111, 8'sb00000010, 8'sb00010000, 8'sb00000000, 8'sb00000100, 8'sb00001011, 8'sb00001110, 8'sb00001110, 8'sb00001001, 8'sb00010101, 8'sb00001111, 8'sb00010011, 8'sb00011010, 8'sb00010100, 8'sb00010001, 8'sb00001010, 8'sb00010001, 8'sb00001001, 8'sb00001011, 8'sb00001111, 8'sb00001110, 8'sb00001111, 8'sb00010011, 8'sb00011011, 8'sb00011110, 8'sb00100101, 8'sb00100100, 8'sb00100101, 8'sb00011101, 8'sb00010001, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00001100, 8'sb00010000, 8'sb00001101, 8'sb00010000, 8'sb00010010, 8'sb00010011, 8'sb00001101, 8'sb00001111, 8'sb00001111, 8'sb00010000, 8'sb00001110, 8'sb00001111,
    8'sb00010000, 8'sb00010010, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00010010, 8'sb00001111, 8'sb00001110, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010110, 8'sb00011111, 8'sb00011100, 8'sb00010010, 8'sb00000100, 8'sb00000101, 8'sb00000111, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00001110, 8'sb00010001, 8'sb00011000, 8'sb00011001, 8'sb00100000, 8'sb00100100, 8'sb00011110, 8'sb00001110, 8'sb00001100, 8'sb00000000, 8'sb00000001, 8'sb00010010, 8'sb00001111, 8'sb00001111, 8'sb00001111, 8'sb00010011, 8'sb00001001, 8'sb00000101, 8'sb00010011, 8'sb00100100, 8'sb00011111, 8'sb00011011, 8'sb00001100, 8'sb00011100, 8'sb00010110, 8'sb00010110, 8'sb00010011, 8'sb00010010, 8'sb00001111, 8'sb00010000, 8'sb00001100, 8'sb00000111, 8'sb00000000, 8'sb00011011, 8'sb00101001, 8'sb00010111, 8'sb00010001, 8'sb00011010, 8'sb00011101, 8'sb00010110, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00001111, 8'sb11111111, 8'sb11111001, 8'sb11100101, 8'sb11101111, 8'sb00011111, 8'sb00011000, 8'sb00010100, 8'sb00000101, 8'sb00000011, 8'sb00010100, 8'sb00001110, 8'sb00001101, 8'sb00001110, 8'sb11111001, 8'sb11100010, 8'sb11111010, 8'sb11111101, 8'sb11111001, 8'sb00011000, 8'sb00000101, 8'sb00001011, 8'sb00000101, 8'sb11111001, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00001111, 8'sb00001010, 8'sb00001010, 8'sb00010000, 8'sb00001010, 8'sb00010001, 8'sb00011011, 8'sb00001010, 8'sb00001100, 8'sb00000100, 8'sb00000010, 8'sb00010101, 8'sb00010100, 8'sb00010001, 8'sb00010110, 8'sb00100010, 8'sb00001010, 8'sb00000100, 8'sb11111100, 8'sb00000001, 8'sb00010000, 8'sb00000101, 8'sb00001001, 8'sb00000111, 8'sb00000111, 8'sb00011000, 8'sb00010001, 8'sb00010001, 8'sb00010100, 8'sb00101001, 8'sb00011001, 8'sb00010111, 8'sb00000101, 8'sb00001110, 8'sb00010111, 8'sb00010010, 8'sb00011001, 8'sb00010001, 8'sb00010111, 8'sb00100000, 8'sb00001111, 8'sb00010000, 8'sb00010100, 8'sb00100001, 8'sb00100101, 8'sb00011101, 8'sb00011001, 8'sb00010000, 8'sb00010001, 8'sb00010100, 8'sb00010110, 8'sb00011000, 8'sb00011001, 8'sb00010110, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00010001, 8'sb00010110, 8'sb00011000, 8'sb00010111, 8'sb00000100, 8'sb00001000, 8'sb00001100, 8'sb00010100, 8'sb00010001, 8'sb00010101, 8'sb00010100, 8'sb00010010, 8'sb00001111, 8'sb00010011, 8'sb00010001, 8'sb00001100, 8'sb00001100, 8'sb00001101, 8'sb00010110, 8'sb00001100, 8'sb00001000, 8'sb00000100, 8'sb00000110, 8'sb00001110, 8'sb00010011, 8'sb00010000, 8'sb00001110, 8'sb00001111, 8'sb00001110, 8'sb00010000, 8'sb00001101, 8'sb00001101, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00010001, 8'sb00001110, 8'sb00001110, 8'sb00010001, 8'sb00001110,
    8'sb00010000, 8'sb00001111, 8'sb00001101, 8'sb00001101, 8'sb00001101, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00001011, 8'sb00001011, 8'sb00001010, 8'sb00001011, 8'sb00001110, 8'sb00011000, 8'sb00010111, 8'sb00010010, 8'sb00001101, 8'sb00010000, 8'sb00001101, 8'sb00001110, 8'sb00010000, 8'sb00001111, 8'sb00001001, 8'sb00001101, 8'sb00001001, 8'sb00001101, 8'sb00010100, 8'sb00100101, 8'sb00100011, 8'sb00100000, 8'sb00011011, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00001011, 8'sb00001100, 8'sb00010001, 8'sb00011001, 8'sb11111001, 8'sb11110001, 8'sb11110111, 8'sb11111100, 8'sb00000011, 8'sb00000110, 8'sb00101001, 8'sb00011000, 8'sb00001111, 8'sb00010000, 8'sb00001011, 8'sb00000111, 8'sb00000100, 8'sb00000110, 8'sb11111011, 8'sb11101011, 8'sb11101101, 8'sb00000100, 8'sb11111111, 8'sb00001010, 8'sb00010001, 8'sb00100001, 8'sb00001111, 8'sb00010000, 8'sb00001011, 8'sb11111111, 8'sb11111010, 8'sb00001000, 8'sb00001110, 8'sb11111111, 8'sb00001111, 8'sb00010001, 8'sb00000000, 8'sb00000001, 8'sb00000111, 8'sb00010100, 8'sb00001110, 8'sb00001111, 8'sb00001101, 8'sb00001011, 8'sb00011010, 8'sb00010100, 8'sb00111001, 8'sb00011100, 8'sb11111110, 8'sb11111100, 8'sb00000010, 8'sb00000111, 8'sb00011001, 8'sb00001111, 8'sb00001100, 8'sb00010000, 8'sb00001110, 8'sb00011110, 8'sb00100001, 8'sb00110000, 8'sb00101011, 8'sb00001111, 8'sb00000110, 8'sb00011000, 8'sb00010101, 8'sb00010100, 8'sb00100110, 8'sb00010110, 8'sb00001100, 8'sb00010000, 8'sb00010010, 8'sb00011000, 8'sb00100011, 8'sb00010100, 8'sb00000110, 8'sb00001110, 8'sb00011010, 8'sb00011100, 8'sb00011010, 8'sb00011110, 8'sb00011111, 8'sb00010001, 8'sb00001100, 8'sb00010000, 8'sb00001110, 8'sb00011111, 8'sb00100010, 8'sb00000011, 8'sb00000001, 8'sb00010010, 8'sb00011101, 8'sb00011000, 8'sb00001110, 8'sb00010010, 8'sb00010100, 8'sb00001011, 8'sb00001011, 8'sb00010000, 8'sb00010000, 8'sb00010111, 8'sb00010110, 8'sb00010111, 8'sb00011010, 8'sb00011101, 8'sb00011101, 8'sb00010111, 8'sb00010011, 8'sb00001101, 8'sb00001111, 8'sb00001100, 8'sb00010000, 8'sb00001101, 8'sb00001100, 8'sb00001100, 8'sb00001011, 8'sb00001001, 8'sb00001101, 8'sb00001101, 8'sb00001000, 8'sb00001110, 8'sb00010110, 8'sb00001110, 8'sb00000011, 8'sb00001110, 8'sb00001101, 8'sb00001111, 8'sb00001101, 8'sb00001100, 8'sb11111111, 8'sb11110010, 8'sb11111010, 8'sb11111110, 8'sb00001000, 8'sb00001000, 8'sb00000110, 8'sb00000100, 8'sb00001001, 8'sb00001101, 8'sb00001111, 8'sb00001111, 8'sb00001100, 8'sb00001110, 8'sb00000111, 8'sb00000111, 8'sb00000010, 8'sb11111111, 8'sb11111010, 8'sb11111111, 8'sb00000001, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00001100,
    8'sb00001111, 8'sb00001100, 8'sb00001111, 8'sb00010000, 8'sb00001100, 8'sb00001110, 8'sb00001101, 8'sb00010001, 8'sb00001110, 8'sb00010000, 8'sb00001101, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00001110, 8'sb00001010, 8'sb00001000, 8'sb00001001, 8'sb00001010, 8'sb00000111, 8'sb00001100, 8'sb00010000, 8'sb00010000, 8'sb00010000, 8'sb00010000, 8'sb00001101, 8'sb00001101, 8'sb00001101, 8'sb00001111, 8'sb00010010, 8'sb00001110, 8'sb00010010, 8'sb00010100, 8'sb00001110, 8'sb00000110, 8'sb00010000, 8'sb00001111, 8'sb00001110, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00010110, 8'sb00011000, 8'sb00010001, 8'sb00000011, 8'sb00011010, 8'sb00100010, 8'sb00010001, 8'sb00000101, 8'sb00001100, 8'sb00010001, 8'sb00001111, 8'sb00001100, 8'sb00010100, 8'sb00011111, 8'sb00011001, 8'sb00011000, 8'sb00001110, 8'sb00001000, 8'sb00100100, 8'sb00011100, 8'sb00010010, 8'sb00001101, 8'sb00000100, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00011001, 8'sb00011011, 8'sb00001111, 8'sb00001101, 8'sb11101010, 8'sb00011011, 8'sb00100100, 8'sb00001011, 8'sb00001100, 8'sb00001111, 8'sb00001001, 8'sb00010000, 8'sb00001110, 8'sb00001101, 8'sb00010010, 8'sb11111011, 8'sb11110011, 8'sb11100110, 8'sb11111110, 8'sb00110010, 8'sb00010011, 8'sb00011100, 8'sb00101011, 8'sb00001111, 8'sb00010001, 8'sb00010000, 8'sb00001101, 8'sb00001101, 8'sb00000100, 8'sb11110011, 8'sb11111001, 8'sb00010000, 8'sb00100111, 8'sb00100100, 8'sb00011100, 8'sb00011111, 8'sb00001011, 8'sb11110110, 8'sb00001010, 8'sb00001110, 8'sb00010001, 8'sb00001011, 8'sb00000101, 8'sb00001011, 8'sb00011100, 8'sb00010111, 8'sb00100100, 8'sb00100000, 8'sb00011001, 8'sb00000110, 8'sb00000000, 8'sb11111011, 8'sb00001110, 8'sb00001101, 8'sb00001111, 8'sb00001100, 8'sb11111101, 8'sb00000000, 8'sb00001000, 8'sb00000000, 8'sb00010001, 8'sb00001100, 8'sb00000000, 8'sb00000110, 8'sb00001001, 8'sb00001010, 8'sb00010010, 8'sb00001101, 8'sb00001101, 8'sb00001111, 8'sb00010011, 8'sb00001111, 8'sb00001011, 8'sb00000001, 8'sb00000001, 8'sb00001000, 8'sb00000110, 8'sb00000101, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00001100, 8'sb00010001, 8'sb00010000, 8'sb00010111, 8'sb00011000, 8'sb00001110, 8'sb00001000, 8'sb00001011, 8'sb00001101, 8'sb00000111, 8'sb00001001, 8'sb00010110, 8'sb00010101, 8'sb00010010, 8'sb00001100, 8'sb00001110, 8'sb00001111, 8'sb00010001, 8'sb00010100, 8'sb00001110, 8'sb00000110, 8'sb00001100, 8'sb00001110, 8'sb00001100, 8'sb00010001, 8'sb00010111, 8'sb00010010, 8'sb00010001, 8'sb00001110, 8'sb00001110, 8'sb00001111, 8'sb00010010, 8'sb00001111, 8'sb00010011, 8'sb00010010, 8'sb00010100, 8'sb00010111, 8'sb00001111, 8'sb00001110, 8'sb00001111, 8'sb00010000, 8'sb00010001, 8'sb00001100,
    8'sb00010000, 8'sb00001101, 8'sb00001110, 8'sb00001101, 8'sb00001111, 8'sb00001100, 8'sb00001101, 8'sb00001101, 8'sb00010000, 8'sb00001111, 8'sb00001100, 8'sb00001111, 8'sb00010000, 8'sb00001011, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00010111, 8'sb00011100, 8'sb00100010, 8'sb00100010, 8'sb00011010, 8'sb00011000, 8'sb00010011, 8'sb00010100, 8'sb00001111, 8'sb00010000, 8'sb00001110, 8'sb00001111, 8'sb00010001, 8'sb00010011, 8'sb00010001, 8'sb00001010, 8'sb00010100, 8'sb00010111, 8'sb00001010, 8'sb00000101, 8'sb00010011, 8'sb00001111, 8'sb00010000, 8'sb00001100, 8'sb00001111, 8'sb00001110, 8'sb00001111, 8'sb00000000, 8'sb00000111, 8'sb00000000, 8'sb00001001, 8'sb00101000, 8'sb00011110, 8'sb11111000, 8'sb00000100, 8'sb11111000, 8'sb00000111, 8'sb00001101, 8'sb00001011, 8'sb00001100, 8'sb00001111, 8'sb00010001, 8'sb00001101, 8'sb11111111, 8'sb00000010, 8'sb00110001, 8'sb00000011, 8'sb11111011, 8'sb00001111, 8'sb11110010, 8'sb11110100, 8'sb00001110, 8'sb00001100, 8'sb00010001, 8'sb00010010, 8'sb00010010, 8'sb11111110, 8'sb11111000, 8'sb11101111, 8'sb01000001, 8'sb00000111, 8'sb00001011, 8'sb00001001, 8'sb00001010, 8'sb00000110, 8'sb00001110, 8'sb00001100, 8'sb00010000, 8'sb00010100, 8'sb00000101, 8'sb00010011, 8'sb00000110, 8'sb11110010, 8'sb00111000, 8'sb00010100, 8'sb00010101, 8'sb00001010, 8'sb00011110, 8'sb00010101, 8'sb00001111, 8'sb00001100, 8'sb00010010, 8'sb00000101, 8'sb00010001, 8'sb00001100, 8'sb00000111, 8'sb00001111, 8'sb00100111, 8'sb00010101, 8'sb00010000, 8'sb00010110, 8'sb00001101, 8'sb00010010, 8'sb00001100, 8'sb00001111, 8'sb00010011, 8'sb00001011, 8'sb00011010, 8'sb00010001, 8'sb00010000, 8'sb00010110, 8'sb00011110, 8'sb00010001, 8'sb00010000, 8'sb00001110, 8'sb00000110, 8'sb00001100, 8'sb00001101, 8'sb00001101, 8'sb00010010, 8'sb00001010, 8'sb00000100, 8'sb00001011, 8'sb00001100, 8'sb00010100, 8'sb00010111, 8'sb00010110, 8'sb00010101, 8'sb00001110, 8'sb00001010, 8'sb00001010, 8'sb00001101, 8'sb00001100, 8'sb00010010, 8'sb00010010, 8'sb00010011, 8'sb00000101, 8'sb00000011, 8'sb00010111, 8'sb00011111, 8'sb00010110, 8'sb00010000, 8'sb00000001, 8'sb11111110, 8'sb00001100, 8'sb00001110, 8'sb00001101, 8'sb00010000, 8'sb00010001, 8'sb00000110, 8'sb11111111, 8'sb11111111, 8'sb00000010, 8'sb00010010, 8'sb00001111, 8'sb00001001, 8'sb00001010, 8'sb00001100, 8'sb00001111, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00010000, 8'sb00010111, 8'sb00010100, 8'sb00011001, 8'sb00001001, 8'sb00001100, 8'sb00010100, 8'sb00011101, 8'sb00100001, 8'sb00010010, 8'sb00001101, 8'sb00001110, 8'sb00001101, 8'sb00001111, 8'sb00001111, 8'sb00010001, 8'sb00011000, 8'sb00011000, 8'sb00010111, 8'sb00011000, 8'sb00010100, 8'sb00010000, 8'sb00010000, 8'sb00010000, 8'sb00001101, 8'sb00001111,
    8'sb00010011, 8'sb00010001, 8'sb00010011, 8'sb00010011, 8'sb00010001, 8'sb00010010, 8'sb00010100, 8'sb00010101, 8'sb00010011, 8'sb00010010, 8'sb00010001, 8'sb00010001, 8'sb00010011, 8'sb00010010, 8'sb00010000, 8'sb00010010, 8'sb00010000, 8'sb00010100, 8'sb00010011, 8'sb00010110, 8'sb00011000, 8'sb00011001, 8'sb00010100, 8'sb00010111, 8'sb00010110, 8'sb00010101, 8'sb00010010, 8'sb00010100, 8'sb00010100, 8'sb00010010, 8'sb00010001, 8'sb00001110, 8'sb00000100, 8'sb11111111, 8'sb00000001, 8'sb00000010, 8'sb00000101, 8'sb00011011, 8'sb00010110, 8'sb00011101, 8'sb00010001, 8'sb00010000, 8'sb00010010, 8'sb00001110, 8'sb00001011, 8'sb11111010, 8'sb11110001, 8'sb00000110, 8'sb00001011, 8'sb00010001, 8'sb00000101, 8'sb00010001, 8'sb00000100, 8'sb00001000, 8'sb00001110, 8'sb00010000, 8'sb00010011, 8'sb00001111, 8'sb11111010, 8'sb11101100, 8'sb00000101, 8'sb00001110, 8'sb00001110, 8'sb00001001, 8'sb00001010, 8'sb11111011, 8'sb11110100, 8'sb00000000, 8'sb00001010, 8'sb00010001, 8'sb00010000, 8'sb00001011, 8'sb11111001, 8'sb00001100, 8'sb00011101, 8'sb00011111, 8'sb00011010, 8'sb00001110, 8'sb11110110, 8'sb00000000, 8'sb00001000, 8'sb00010100, 8'sb00001000, 8'sb00010000, 8'sb00010000, 8'sb00001100, 8'sb00010001, 8'sb00101000, 8'sb00011110, 8'sb00001110, 8'sb00010011, 8'sb00011010, 8'sb00010010, 8'sb00010100, 8'sb00010101, 8'sb00101100, 8'sb00011010, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00001110, 8'sb00100011, 8'sb00011001, 8'sb00001100, 8'sb00001000, 8'sb00011110, 8'sb00011000, 8'sb11111111, 8'sb00001110, 8'sb00010011, 8'sb00001110, 8'sb00001101, 8'sb00010100, 8'sb00001101, 8'sb11111011, 8'sb00001010, 8'sb00011100, 8'sb00100010, 8'sb00010011, 8'sb00011111, 8'sb00000010, 8'sb00000101, 8'sb00000001, 8'sb00000110, 8'sb00001000, 8'sb00010001, 8'sb00010011, 8'sb00001101, 8'sb11111101, 8'sb11111000, 8'sb11111110, 8'sb00001101, 8'sb00011000, 8'sb00001111, 8'sb00000101, 8'sb00000101, 8'sb00001111, 8'sb00001100, 8'sb00000100, 8'sb00010010, 8'sb00001111, 8'sb00010001, 8'sb00000100, 8'sb00001000, 8'sb00001110, 8'sb00011000, 8'sb00011001, 8'sb00011010, 8'sb00010100, 8'sb00001010, 8'sb00001101, 8'sb00001001, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00010000, 8'sb00001110, 8'sb00000100, 8'sb00011010, 8'sb00001111, 8'sb00010001, 8'sb00001101, 8'sb00010111, 8'sb00000110, 8'sb00000111, 8'sb00001101, 8'sb00010001, 8'sb00010000, 8'sb00010010, 8'sb00010100, 8'sb00010101, 8'sb00010000, 8'sb00010001, 8'sb00001010, 8'sb00000100, 8'sb00000101, 8'sb00001101, 8'sb00001110, 8'sb00010101, 8'sb00010110, 8'sb00010010, 8'sb00010001, 8'sb00010011, 8'sb00010100, 8'sb00010001, 8'sb00010101, 8'sb00010011, 8'sb00010100, 8'sb00010101, 8'sb00010101, 8'sb00010001, 8'sb00001111, 8'sb00010001, 8'sb00010011, 8'sb00010001, 8'sb00010100,
    8'sb00001010, 8'sb00001101, 8'sb00001011, 8'sb00001001, 8'sb00001011, 8'sb00001010, 8'sb00001011, 8'sb00001011, 8'sb00001000, 8'sb00001011, 8'sb00001100, 8'sb00001010, 8'sb00001011, 8'sb00001100, 8'sb00001001, 8'sb00001101, 8'sb00001000, 8'sb00001010, 8'sb00001100, 8'sb00001010, 8'sb11111111, 8'sb00000000, 8'sb00001011, 8'sb00010001, 8'sb00001110, 8'sb00001011, 8'sb00001001, 8'sb00001011, 8'sb00001001, 8'sb00001001, 8'sb00001000, 8'sb00000101, 8'sb00001010, 8'sb00001000, 8'sb00001100, 8'sb00001011, 8'sb00010101, 8'sb00011011, 8'sb00011001, 8'sb00010110, 8'sb00001110, 8'sb00001011, 8'sb00001010, 8'sb00001010, 8'sb00000100, 8'sb00010000, 8'sb00010000, 8'sb00001101, 8'sb00010000, 8'sb00001110, 8'sb00010111, 8'sb00010011, 8'sb00101111, 8'sb00101111, 8'sb00010100, 8'sb00001110, 8'sb00001010, 8'sb00001000, 8'sb00000001, 8'sb00001001, 8'sb00011000, 8'sb00011101, 8'sb00010010, 8'sb11110011, 8'sb11110010, 8'sb00010000, 8'sb00111111, 8'sb00110100, 8'sb00011001, 8'sb00001011, 8'sb00001001, 8'sb00001000, 8'sb00010000, 8'sb00100000, 8'sb00100100, 8'sb00000101, 8'sb00000100, 8'sb11101001, 8'sb00001011, 8'sb00101100, 8'sb00110011, 8'sb00011100, 8'sb00010010, 8'sb00001010, 8'sb00001101, 8'sb00001100, 8'sb00011000, 8'sb00011010, 8'sb00001000, 8'sb00010001, 8'sb11111101, 8'sb00000011, 8'sb00011101, 8'sb00101001, 8'sb00100000, 8'sb00010000, 8'sb00001010, 8'sb00001011, 8'sb00001000, 8'sb00001101, 8'sb00010000, 8'sb00010000, 8'sb00001001, 8'sb00010100, 8'sb00001010, 8'sb00001111, 8'sb00011100, 8'sb00011000, 8'sb00001000, 8'sb00001100, 8'sb00010000, 8'sb00001011, 8'sb00001000, 8'sb00001010, 8'sb00010010, 8'sb00010010, 8'sb00001001, 8'sb00001001, 8'sb00010011, 8'sb00011001, 8'sb00011101, 8'sb00001101, 8'sb00001000, 8'sb11111111, 8'sb00001111, 8'sb00001001, 8'sb00001010, 8'sb00000111, 8'sb00010011, 8'sb00010010, 8'sb00010011, 8'sb00010011, 8'sb00001011, 8'sb00001111, 8'sb00000101, 8'sb00001000, 8'sb00000100, 8'sb00000100, 8'sb00001110, 8'sb00001100, 8'sb00001001, 8'sb00001001, 8'sb00010100, 8'sb00010111, 8'sb00010100, 8'sb00010100, 8'sb00011010, 8'sb00001110, 8'sb00001100, 8'sb00001111, 8'sb00010101, 8'sb00011011, 8'sb00001101, 8'sb00001011, 8'sb00001011, 8'sb00000110, 8'sb00001000, 8'sb00010011, 8'sb00001100, 8'sb00001010, 8'sb00010010, 8'sb00011000, 8'sb00001001, 8'sb00000001, 8'sb00010110, 8'sb00010000, 8'sb00001101, 8'sb00001010, 8'sb00001001, 8'sb00001001, 8'sb00000101, 8'sb00000100, 8'sb00000101, 8'sb00001111, 8'sb00001111, 8'sb00010000, 8'sb00001110, 8'sb00010010, 8'sb00010000, 8'sb00001010, 8'sb00001000, 8'sb00001011, 8'sb00001000, 8'sb00001100, 8'sb00001000, 8'sb00001010, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00001110, 8'sb00001011, 8'sb00001010, 8'sb00001010, 8'sb00001101, 8'sb00001010, 8'sb00001010,
    8'sb00001110, 8'sb00001111, 8'sb00001111, 8'sb00001011, 8'sb00001011, 8'sb00001110, 8'sb00001111, 8'sb00001111, 8'sb00001111, 8'sb00001011, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00001100, 8'sb00001110, 8'sb00001011, 8'sb00001101, 8'sb00010011, 8'sb00010100, 8'sb00010111, 8'sb00011011, 8'sb00011000, 8'sb00001100, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00001001, 8'sb00000110, 8'sb00001110, 8'sb00010000, 8'sb00010100, 8'sb00011011, 8'sb00010100, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00010010, 8'sb00001110, 8'sb00001100, 8'sb00001100, 8'sb00001011, 8'sb11111101, 8'sb00001001, 8'sb00001111, 8'sb00000111, 8'sb00000011, 8'sb00010111, 8'sb00011101, 8'sb00000101, 8'sb00001001, 8'sb00001110, 8'sb00011100, 8'sb00001100, 8'sb00001111, 8'sb00001010, 8'sb11111100, 8'sb11111110, 8'sb00000000, 8'sb00001011, 8'sb00001111, 8'sb00010101, 8'sb00000100, 8'sb00000110, 8'sb00001001, 8'sb00100100, 8'sb00101111, 8'sb00001100, 8'sb00001011, 8'sb00001011, 8'sb00010000, 8'sb00100000, 8'sb00101000, 8'sb00101001, 8'sb00110010, 8'sb00001101, 8'sb11110000, 8'sb00000011, 8'sb00010111, 8'sb00100110, 8'sb00011100, 8'sb00001111, 8'sb00001100, 8'sb00001101, 8'sb00011100, 8'sb00101110, 8'sb00100100, 8'sb00011010, 8'sb00011110, 8'sb00011010, 8'sb00001000, 8'sb00001001, 8'sb00010100, 8'sb00011001, 8'sb00001110, 8'sb00001110, 8'sb00001100, 8'sb00001010, 8'sb00001010, 8'sb00000111, 8'sb00010001, 8'sb00001110, 8'sb00010110, 8'sb11111111, 8'sb00000111, 8'sb00000001, 8'sb00000001, 8'sb00010110, 8'sb00001100, 8'sb00001100, 8'sb00001100, 8'sb00000110, 8'sb00000110, 8'sb00001011, 8'sb00010110, 8'sb00011010, 8'sb00001000, 8'sb11111101, 8'sb00000011, 8'sb11111111, 8'sb00000101, 8'sb00010000, 8'sb00001110, 8'sb00001110, 8'sb00001011, 8'sb00001001, 8'sb00000111, 8'sb00001101, 8'sb00010011, 8'sb00100111, 8'sb00010011, 8'sb11111110, 8'sb00010011, 8'sb00010100, 8'sb00010100, 8'sb00010110, 8'sb00001010, 8'sb00001110, 8'sb00001101, 8'sb00001000, 8'sb00000110, 8'sb00000110, 8'sb00001110, 8'sb00010111, 8'sb00011010, 8'sb00000010, 8'sb00000111, 8'sb00000111, 8'sb00001100, 8'sb00010111, 8'sb00001101, 8'sb00001011, 8'sb00001011, 8'sb00001010, 8'sb00000111, 8'sb00000101, 8'sb00010001, 8'sb00011011, 8'sb00100010, 8'sb00001011, 8'sb00000110, 8'sb00000000, 8'sb00001011, 8'sb00001101, 8'sb00001001, 8'sb00001101, 8'sb00001010, 8'sb00001101, 8'sb00000111, 8'sb00001001, 8'sb00010100, 8'sb00011001, 8'sb00011101, 8'sb00010010, 8'sb00010110, 8'sb00010010, 8'sb00001101, 8'sb00001010, 8'sb00001011, 8'sb00001111, 8'sb00001011, 8'sb00001110, 8'sb00001100, 8'sb00001011, 8'sb00001101, 8'sb00010001, 8'sb00010101, 8'sb00010001, 8'sb00001111, 8'sb00001101, 8'sb00001101, 8'sb00001101, 8'sb00001100, 8'sb00001110,
    8'sb00010011, 8'sb00010011, 8'sb00010011, 8'sb00001110, 8'sb00010000, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00010001, 8'sb00010001, 8'sb00010001, 8'sb00010000, 8'sb00010000, 8'sb00010010, 8'sb00010011, 8'sb00010000, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00010001, 8'sb00010011, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00001101, 8'sb00001101, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00010001, 8'sb00010001, 8'sb00001111, 8'sb00001010, 8'sb00001100, 8'sb00010011, 8'sb00011000, 8'sb00100100, 8'sb00010110, 8'sb00010010, 8'sb00000100, 8'sb00010011, 8'sb00010100, 8'sb00010000, 8'sb00010010, 8'sb00010001, 8'sb00001001, 8'sb00000100, 8'sb00001110, 8'sb00000110, 8'sb00001100, 8'sb00011110, 8'sb00011101, 8'sb00010110, 8'sb00001110, 8'sb00000111, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00010001, 8'sb00010100, 8'sb00010110, 8'sb00001111, 8'sb00010010, 8'sb11111111, 8'sb00001010, 8'sb00110101, 8'sb00011000, 8'sb00011010, 8'sb11110011, 8'sb00001100, 8'sb00010000, 8'sb00001011, 8'sb00001110, 8'sb00001111, 8'sb00010111, 8'sb00001010, 8'sb00000111, 8'sb11011000, 8'sb00101010, 8'sb00101111, 8'sb00011110, 8'sb00011111, 8'sb11110011, 8'sb00001010, 8'sb00001111, 8'sb00001111, 8'sb00001000, 8'sb00001011, 8'sb00001000, 8'sb11111110, 8'sb00000001, 8'sb00000111, 8'sb00100110, 8'sb00100100, 8'sb00100111, 8'sb01000001, 8'sb00110010, 8'sb00001110, 8'sb00010010, 8'sb00001110, 8'sb00010101, 8'sb00011101, 8'sb00000010, 8'sb00001000, 8'sb00001111, 8'sb00010101, 8'sb00010100, 8'sb00010010, 8'sb00001001, 8'sb00001111, 8'sb00011010, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00010110, 8'sb00011101, 8'sb00001010, 8'sb00010111, 8'sb00001101, 8'sb00011000, 8'sb00001000, 8'sb00001011, 8'sb00001010, 8'sb00001011, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00000100, 8'sb00000100, 8'sb00010100, 8'sb00010100, 8'sb00001100, 8'sb00001001, 8'sb00001000, 8'sb00000111, 8'sb00000000, 8'sb11111110, 8'sb00001110, 8'sb00010010, 8'sb00001111, 8'sb00010010, 8'sb00001101, 8'sb00011100, 8'sb00001101, 8'sb00010001, 8'sb00010010, 8'sb00010011, 8'sb00000100, 8'sb00000110, 8'sb00000010, 8'sb11111111, 8'sb00001110, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00001000, 8'sb00010101, 8'sb00001000, 8'sb00001100, 8'sb00010110, 8'sb00001110, 8'sb00000100, 8'sb00001011, 8'sb00001011, 8'sb00001110, 8'sb00010100, 8'sb00010000, 8'sb00010010, 8'sb00001111, 8'sb00001101, 8'sb00001011, 8'sb00001001, 8'sb00010001, 8'sb00010001, 8'sb00010011, 8'sb00010000, 8'sb00010001, 8'sb00001100, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00010001, 8'sb00010001, 8'sb00001110, 8'sb00010010, 8'sb00010001, 8'sb00010000, 8'sb00001110, 8'sb00001011, 8'sb00001110, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00010000,
    8'sb00010001, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00001100, 8'sb00001011, 8'sb00001010, 8'sb00001011, 8'sb00001011, 8'sb00001001, 8'sb00001110, 8'sb00010010, 8'sb00010001, 8'sb00001101, 8'sb00001101, 8'sb00010000, 8'sb00001101, 8'sb00001010, 8'sb00000000, 8'sb00000010, 8'sb00001001, 8'sb00001001, 8'sb00000110, 8'sb00001111, 8'sb00010000, 8'sb00010111, 8'sb00100010, 8'sb00010010, 8'sb00010001, 8'sb00001110, 8'sb00001101, 8'sb00000001, 8'sb00000110, 8'sb00010100, 8'sb00011011, 8'sb00011010, 8'sb00001000, 8'sb00001001, 8'sb00010000, 8'sb00001101, 8'sb00011001, 8'sb00011000, 8'sb00001110, 8'sb00010000, 8'sb00001100, 8'sb00000000, 8'sb00001011, 8'sb00010001, 8'sb00100000, 8'sb00001100, 8'sb00001110, 8'sb00010110, 8'sb00010101, 8'sb00010001, 8'sb00001110, 8'sb00011011, 8'sb00001111, 8'sb00010000, 8'sb00001101, 8'sb00010001, 8'sb00011000, 8'sb00010111, 8'sb00101110, 8'sb00001001, 8'sb11110001, 8'sb00010110, 8'sb00000100, 8'sb00000100, 8'sb00000101, 8'sb00001110, 8'sb00001111, 8'sb00001111, 8'sb00010001, 8'sb00011110, 8'sb00101100, 8'sb00100000, 8'sb00100001, 8'sb11111111, 8'sb11110100, 8'sb00010110, 8'sb00011100, 8'sb00010110, 8'sb00010110, 8'sb00001011, 8'sb00001101, 8'sb00010001, 8'sb00010000, 8'sb00100000, 8'sb00100011, 8'sb00010111, 8'sb00010001, 8'sb11111111, 8'sb11101000, 8'sb00010111, 8'sb00001101, 8'sb00010001, 8'sb00010111, 8'sb00010010, 8'sb00001101, 8'sb00001101, 8'sb00001010, 8'sb00010111, 8'sb00010110, 8'sb00001101, 8'sb00001100, 8'sb11110000, 8'sb11111101, 8'sb00011100, 8'sb00010010, 8'sb00010100, 8'sb00000010, 8'sb00001100, 8'sb00001101, 8'sb00001111, 8'sb00000111, 8'sb00001111, 8'sb00001111, 8'sb00001001, 8'sb00000000, 8'sb11101100, 8'sb00010101, 8'sb00001110, 8'sb00001110, 8'sb00000110, 8'sb11111110, 8'sb00001010, 8'sb00001100, 8'sb00010001, 8'sb00001100, 8'sb00010110, 8'sb00001111, 8'sb11111111, 8'sb11111100, 8'sb00010100, 8'sb00010011, 8'sb00001110, 8'sb00001010, 8'sb00000010, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010001, 8'sb00001011, 8'sb00001001, 8'sb00000100, 8'sb00000100, 8'sb00000101, 8'sb00011001, 8'sb00010011, 8'sb00010011, 8'sb00010001, 8'sb00010100, 8'sb00010100, 8'sb00001111, 8'sb00001101, 8'sb00010001, 8'sb00001100, 8'sb00001110, 8'sb00001000, 8'sb00001011, 8'sb00001101, 8'sb00001111, 8'sb00010001, 8'sb00010100, 8'sb00010100, 8'sb00010111, 8'sb00010001, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00001101, 8'sb00010001, 8'sb00010001, 8'sb00010010, 8'sb00010101, 8'sb00010011, 8'sb00010011, 8'sb00010011, 8'sb00010011, 8'sb00001110, 8'sb00010010, 8'sb00010000, 8'sb00010001,
    8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00001011, 8'sb00001010, 8'sb00001010, 8'sb00001100, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00001110, 8'sb00001011, 8'sb00001010, 8'sb00001110, 8'sb00001100, 8'sb00001110, 8'sb00001100, 8'sb00001111, 8'sb00001101, 8'sb00001100, 8'sb00010010, 8'sb00001111, 8'sb00001100, 8'sb00000110, 8'sb00001000, 8'sb00001100, 8'sb00001010, 8'sb00001010, 8'sb00001101, 8'sb00001110, 8'sb00001101, 8'sb00001110, 8'sb00010010, 8'sb00010001, 8'sb00001001, 8'sb00000111, 8'sb11110111, 8'sb00001100, 8'sb11111111, 8'sb11111101, 8'sb00001100, 8'sb00001100, 8'sb00001011, 8'sb00001101, 8'sb00001010, 8'sb00001001, 8'sb00010010, 8'sb00011000, 8'sb00101101, 8'sb00100100, 8'sb00100101, 8'sb00100101, 8'sb00100101, 8'sb11111101, 8'sb00000011, 8'sb00001010, 8'sb00001101, 8'sb00001010, 8'sb00000001, 8'sb00001001, 8'sb00010101, 8'sb00010100, 8'sb00100011, 8'sb00110111, 8'sb00101010, 8'sb00011000, 8'sb00010000, 8'sb00011011, 8'sb00001110, 8'sb00001011, 8'sb00001101, 8'sb00001111, 8'sb00001100, 8'sb00011010, 8'sb00010111, 8'sb00011110, 8'sb00101001, 8'sb00011110, 8'sb00010110, 8'sb00011001, 8'sb00011011, 8'sb00100011, 8'sb00011000, 8'sb00001011, 8'sb00001100, 8'sb00010011, 8'sb00011111, 8'sb00010100, 8'sb00010101, 8'sb00000110, 8'sb11101010, 8'sb00000110, 8'sb00001110, 8'sb00010010, 8'sb00010000, 8'sb00001111, 8'sb00000101, 8'sb00001101, 8'sb00001110, 8'sb00001110, 8'sb00010001, 8'sb00001011, 8'sb00000010, 8'sb00000001, 8'sb11110101, 8'sb11110111, 8'sb00000100, 8'sb11111101, 8'sb00001101, 8'sb11111101, 8'sb00000100, 8'sb00001100, 8'sb00001100, 8'sb00001101, 8'sb00001100, 8'sb11111101, 8'sb00000011, 8'sb00011000, 8'sb11111100, 8'sb11101110, 8'sb00000001, 8'sb00000110, 8'sb11111010, 8'sb11111100, 8'sb00000101, 8'sb00001010, 8'sb00001110, 8'sb00000111, 8'sb00001100, 8'sb00001100, 8'sb00010010, 8'sb00001100, 8'sb11111100, 8'sb00001001, 8'sb00001001, 8'sb00011001, 8'sb00010110, 8'sb00001111, 8'sb00000111, 8'sb00001101, 8'sb00001010, 8'sb00001011, 8'sb00010011, 8'sb00010101, 8'sb00010100, 8'sb11111010, 8'sb00000010, 8'sb00001001, 8'sb00001000, 8'sb00010001, 8'sb00010101, 8'sb00010110, 8'sb00001110, 8'sb00001010, 8'sb00001101, 8'sb00001011, 8'sb00001111, 8'sb00011010, 8'sb00011110, 8'sb00001100, 8'sb00001000, 8'sb00000000, 8'sb11111100, 8'sb11110111, 8'sb00000011, 8'sb00011010, 8'sb00001110, 8'sb00001011, 8'sb00001011, 8'sb00001011, 8'sb00010001, 8'sb00011110, 8'sb00100010, 8'sb00011101, 8'sb00011111, 8'sb00100010, 8'sb00100110, 8'sb00100010, 8'sb00010101, 8'sb00010110, 8'sb00001111, 8'sb00001011, 8'sb00001101, 8'sb00001110, 8'sb00001111, 8'sb00010100, 8'sb00011000, 8'sb00011011, 8'sb00100000, 8'sb00100100, 8'sb00100001, 8'sb00011010, 8'sb00010000, 8'sb00001111, 8'sb00001100, 8'sb00001100,
    8'sb00010100, 8'sb00010000, 8'sb00001111, 8'sb00010011, 8'sb00010011, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00010010, 8'sb00010000, 8'sb00010000, 8'sb00010001, 8'sb00010011, 8'sb00010001, 8'sb00010100, 8'sb00010100, 8'sb00010010, 8'sb00010000, 8'sb00001111, 8'sb00001100, 8'sb00001001, 8'sb00001001, 8'sb00001110, 8'sb00010101, 8'sb00010100, 8'sb00010111, 8'sb00010001, 8'sb00010001, 8'sb00010010, 8'sb00010010, 8'sb00010100, 8'sb00010011, 8'sb00001010, 8'sb00000010, 8'sb00000110, 8'sb00010000, 8'sb00000111, 8'sb00001101, 8'sb00011010, 8'sb00011011, 8'sb00001110, 8'sb00010010, 8'sb00010011, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00000100, 8'sb11111111, 8'sb11110010, 8'sb11100111, 8'sb11101011, 8'sb00000010, 8'sb00001101, 8'sb00010100, 8'sb00001100, 8'sb00001110, 8'sb00001111, 8'sb00010000, 8'sb00010001, 8'sb00000011, 8'sb11111000, 8'sb11101101, 8'sb11110101, 8'sb00000000, 8'sb00010010, 8'sb00000100, 8'sb00000110, 8'sb11111000, 8'sb11111000, 8'sb00001011, 8'sb00010011, 8'sb00010010, 8'sb00001110, 8'sb00010001, 8'sb00100001, 8'sb00110110, 8'sb00111111, 8'sb00011010, 8'sb00000101, 8'sb00000110, 8'sb00010011, 8'sb00000010, 8'sb11111101, 8'sb00001111, 8'sb00010000, 8'sb00010000, 8'sb00011011, 8'sb00100111, 8'sb00101010, 8'sb00011010, 8'sb00001011, 8'sb00010001, 8'sb00010011, 8'sb00001101, 8'sb00001111, 8'sb00011011, 8'sb00010011, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00011100, 8'sb00010110, 8'sb00001100, 8'sb00000111, 8'sb00011001, 8'sb00010110, 8'sb00001111, 8'sb00010010, 8'sb00010110, 8'sb00011010, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00001100, 8'sb11111011, 8'sb00001110, 8'sb00011011, 8'sb00010111, 8'sb00011010, 8'sb00010001, 8'sb00001000, 8'sb00010010, 8'sb00010011, 8'sb00000100, 8'sb11111111, 8'sb00001111, 8'sb00010010, 8'sb00001101, 8'sb11110011, 8'sb11101010, 8'sb00010010, 8'sb00010111, 8'sb00011100, 8'sb00001111, 8'sb00001100, 8'sb00010010, 8'sb00001100, 8'sb00000000, 8'sb00000000, 8'sb00010001, 8'sb00010010, 8'sb00001100, 8'sb00000000, 8'sb11111101, 8'sb00000001, 8'sb00001010, 8'sb00010011, 8'sb00011000, 8'sb00010110, 8'sb00010100, 8'sb00000010, 8'sb11111111, 8'sb00001101, 8'sb00010011, 8'sb00001111, 8'sb00010001, 8'sb00010100, 8'sb00010100, 8'sb00001111, 8'sb00001111, 8'sb00010100, 8'sb00011001, 8'sb00010111, 8'sb00011000, 8'sb00001000, 8'sb00000110, 8'sb00001101, 8'sb00010001, 8'sb00010010, 8'sb00010000, 8'sb00010010, 8'sb00001111, 8'sb00001100, 8'sb00010100, 8'sb00001010, 8'sb00001001, 8'sb00000110, 8'sb00001001, 8'sb00001001, 8'sb00001110, 8'sb00001101, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00010000, 8'sb00001111, 8'sb00001010, 8'sb00000101, 8'sb00001000, 8'sb00001100, 8'sb00001100, 8'sb00010001, 8'sb00010010, 8'sb00001111,
    8'sb00010011, 8'sb00010000, 8'sb00010000, 8'sb00010001, 8'sb00010000, 8'sb00010010, 8'sb00010000, 8'sb00010011, 8'sb00001111, 8'sb00010001, 8'sb00010010, 8'sb00010010, 8'sb00010011, 8'sb00010001, 8'sb00010010, 8'sb00001111, 8'sb00010001, 8'sb00010010, 8'sb00010001, 8'sb00010010, 8'sb00010101, 8'sb00010110, 8'sb00011010, 8'sb00010011, 8'sb00010010, 8'sb00010100, 8'sb00010001, 8'sb00010010, 8'sb00010100, 8'sb00010011, 8'sb00010100, 8'sb00001110, 8'sb00001111, 8'sb00001011, 8'sb00001001, 8'sb00001000, 8'sb11111110, 8'sb00000101, 8'sb00010000, 8'sb00010011, 8'sb00001010, 8'sb00010011, 8'sb00010000, 8'sb00001110, 8'sb00001001, 8'sb11111001, 8'sb11110101, 8'sb11111110, 8'sb11111100, 8'sb00001010, 8'sb00000101, 8'sb00000100, 8'sb00001001, 8'sb00000110, 8'sb00000110, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb11111010, 8'sb11110110, 8'sb11110101, 8'sb00000010, 8'sb00010000, 8'sb00010001, 8'sb11111011, 8'sb00000101, 8'sb00001000, 8'sb11111001, 8'sb11111110, 8'sb00010000, 8'sb00010011, 8'sb00001011, 8'sb00001010, 8'sb00001001, 8'sb00001011, 8'sb00000011, 8'sb11110101, 8'sb00000011, 8'sb00001011, 8'sb00001001, 8'sb00000111, 8'sb11110111, 8'sb11111111, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00011110, 8'sb00100011, 8'sb00011010, 8'sb00010101, 8'sb00110000, 8'sb00101101, 8'sb00010001, 8'sb00100001, 8'sb00100101, 8'sb00010000, 8'sb00001100, 8'sb00010000, 8'sb00010001, 8'sb00010010, 8'sb00100010, 8'sb00100111, 8'sb00100000, 8'sb00011011, 8'sb00100100, 8'sb00011110, 8'sb00011001, 8'sb00010011, 8'sb00010101, 8'sb00001001, 8'sb00010010, 8'sb00010011, 8'sb00010011, 8'sb00010010, 8'sb00011010, 8'sb00011100, 8'sb00001001, 8'sb00010100, 8'sb00011011, 8'sb00100010, 8'sb00010111, 8'sb00001110, 8'sb00001101, 8'sb00001001, 8'sb00001110, 8'sb00010010, 8'sb00010011, 8'sb00001111, 8'sb00000101, 8'sb00001000, 8'sb00011100, 8'sb00011110, 8'sb00100100, 8'sb00101011, 8'sb00011011, 8'sb00010010, 8'sb00001011, 8'sb00000111, 8'sb00010101, 8'sb00010100, 8'sb00010000, 8'sb00010001, 8'sb00000010, 8'sb11101010, 8'sb11101111, 8'sb00000001, 8'sb00001000, 8'sb00000111, 8'sb00000110, 8'sb00001100, 8'sb00000000, 8'sb00001000, 8'sb00010010, 8'sb00010010, 8'sb00010010, 8'sb00010001, 8'sb00001100, 8'sb00000000, 8'sb11110111, 8'sb11100101, 8'sb11100100, 8'sb11101101, 8'sb11101111, 8'sb11111100, 8'sb00000110, 8'sb00001111, 8'sb00010011, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00001111, 8'sb00001001, 8'sb11111111, 8'sb11111100, 8'sb00010000, 8'sb00010000, 8'sb00011110, 8'sb00010100, 8'sb00010011, 8'sb00010011, 8'sb00010010, 8'sb00010100, 8'sb00010001, 8'sb00010010, 8'sb00001101, 8'sb00001110, 8'sb00010100, 8'sb00010101, 8'sb00010000, 8'sb00001110, 8'sb00010011, 8'sb00010010, 8'sb00010001, 8'sb00010000,
    8'sb00001100, 8'sb00001101, 8'sb00001101, 8'sb00001101, 8'sb00001011, 8'sb00001011, 8'sb00001110, 8'sb00001100, 8'sb00001010, 8'sb00001011, 8'sb00001100, 8'sb00001011, 8'sb00001111, 8'sb00001111, 8'sb00001101, 8'sb00001111, 8'sb00001110, 8'sb00001101, 8'sb00001111, 8'sb00010110, 8'sb00011010, 8'sb00010011, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00001110, 8'sb00001101, 8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00001111, 8'sb00010100, 8'sb00011000, 8'sb00011110, 8'sb00011000, 8'sb00000010, 8'sb00001111, 8'sb00010111, 8'sb00010101, 8'sb00001111, 8'sb00010011, 8'sb00001101, 8'sb00001110, 8'sb00001011, 8'sb00010000, 8'sb00010010, 8'sb00011111, 8'sb00001100, 8'sb00001100, 8'sb00010111, 8'sb00010010, 8'sb00000100, 8'sb00000111, 8'sb00001101, 8'sb00010011, 8'sb00001011, 8'sb00001100, 8'sb00001010, 8'sb00000101, 8'sb00001010, 8'sb00001111, 8'sb00010000, 8'sb00000111, 8'sb00000000, 8'sb11111111, 8'sb00000001, 8'sb00000100, 8'sb00000111, 8'sb00000110, 8'sb00001111, 8'sb00001011, 8'sb00000111, 8'sb00001000, 8'sb00010100, 8'sb00100010, 8'sb00010100, 8'sb11110000, 8'sb11101110, 8'sb00000001, 8'sb00000100, 8'sb00000010, 8'sb11111101, 8'sb00000010, 8'sb00001110, 8'sb00001011, 8'sb00001010, 8'sb00000110, 8'sb00000100, 8'sb00010100, 8'sb00101011, 8'sb00011010, 8'sb00001100, 8'sb00010010, 8'sb00010100, 8'sb00010000, 8'sb00001000, 8'sb00001111, 8'sb00001111, 8'sb00001111, 8'sb00001111, 8'sb00000110, 8'sb00001111, 8'sb00010000, 8'sb00011110, 8'sb00100010, 8'sb00010011, 8'sb00011001, 8'sb00001011, 8'sb00001001, 8'sb00001100, 8'sb00001110, 8'sb00001110, 8'sb00001100, 8'sb00001110, 8'sb00001100, 8'sb00000110, 8'sb00010011, 8'sb00011010, 8'sb00101011, 8'sb00010110, 8'sb00011011, 8'sb00011101, 8'sb00011000, 8'sb00011000, 8'sb00010110, 8'sb00010000, 8'sb00001111, 8'sb00010011, 8'sb00011011, 8'sb00010011, 8'sb11111111, 8'sb00001100, 8'sb00001111, 8'sb00001011, 8'sb00010001, 8'sb00010000, 8'sb00011000, 8'sb00010111, 8'sb00011000, 8'sb00001110, 8'sb00001011, 8'sb00010011, 8'sb00011000, 8'sb00001101, 8'sb00001010, 8'sb11111101, 8'sb00010100, 8'sb00011100, 8'sb00010001, 8'sb00011001, 8'sb00011000, 8'sb00011111, 8'sb00001111, 8'sb00001111, 8'sb00001101, 8'sb00010001, 8'sb00010110, 8'sb00001100, 8'sb00010110, 8'sb00010010, 8'sb00001000, 8'sb00001101, 8'sb00010101, 8'sb00101001, 8'sb00100011, 8'sb00010111, 8'sb00010000, 8'sb00001101, 8'sb00001100, 8'sb00001111, 8'sb00001101, 8'sb00001001, 8'sb00001100, 8'sb00010011, 8'sb00010010, 8'sb00010100, 8'sb00001110, 8'sb00010100, 8'sb00010101, 8'sb00010011, 8'sb00001111, 8'sb00001110, 8'sb00001100, 8'sb00001011, 8'sb00001110, 8'sb00001101, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00001101, 8'sb00000110, 8'sb00000101, 8'sb00001101, 8'sb00001110, 8'sb00001111, 8'sb00001100,
    8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00001101, 8'sb00001101, 8'sb00010001, 8'sb00001101, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00001101, 8'sb00001110, 8'sb00001110, 8'sb00001101, 8'sb00010000, 8'sb00001110, 8'sb00001100, 8'sb00010001, 8'sb00001110, 8'sb00000111, 8'sb00001010, 8'sb00001001, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00001111, 8'sb00001101, 8'sb00001101, 8'sb00001101, 8'sb00001100, 8'sb11111111, 8'sb11111100, 8'sb00000001, 8'sb00000011, 8'sb00010100, 8'sb00011110, 8'sb00010100, 8'sb00010001, 8'sb00001111, 8'sb00001101, 8'sb00001011, 8'sb00010011, 8'sb00011010, 8'sb00100000, 8'sb00010100, 8'sb11111111, 8'sb11110011, 8'sb00000101, 8'sb00001001, 8'sb00011101, 8'sb00100011, 8'sb00010000, 8'sb00001111, 8'sb00001101, 8'sb00001111, 8'sb00001101, 8'sb00010001, 8'sb00010110, 8'sb00101110, 8'sb00000000, 8'sb11100100, 8'sb11110100, 8'sb00000110, 8'sb00001010, 8'sb00100110, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00010100, 8'sb00010101, 8'sb00010010, 8'sb00100010, 8'sb00101010, 8'sb00000001, 8'sb11101110, 8'sb11111000, 8'sb00000011, 8'sb00010110, 8'sb00010010, 8'sb00001100, 8'sb00001100, 8'sb00001111, 8'sb00011000, 8'sb00010001, 8'sb00001110, 8'sb00100011, 8'sb00100001, 8'sb00010010, 8'sb00001010, 8'sb00001101, 8'sb00000110, 8'sb00001100, 8'sb00001101, 8'sb00001110, 8'sb00001110, 8'sb00001000, 8'sb00000111, 8'sb00001110, 8'sb00011100, 8'sb00011100, 8'sb00100101, 8'sb00000100, 8'sb00001100, 8'sb00001001, 8'sb00001000, 8'sb00010000, 8'sb00001110, 8'sb00001101, 8'sb00001100, 8'sb00000010, 8'sb00001010, 8'sb00010011, 8'sb00010101, 8'sb00100101, 8'sb00011011, 8'sb00001101, 8'sb00001001, 8'sb00010000, 8'sb00010001, 8'sb00010011, 8'sb00001101, 8'sb00010000, 8'sb00001101, 8'sb00001111, 8'sb00010001, 8'sb00011000, 8'sb00010100, 8'sb00001110, 8'sb00010010, 8'sb00001110, 8'sb00001110, 8'sb00010100, 8'sb00011000, 8'sb00001101, 8'sb00010000, 8'sb00010001, 8'sb00001001, 8'sb00001000, 8'sb00010011, 8'sb00010100, 8'sb00001011, 8'sb00000100, 8'sb00010101, 8'sb00010100, 8'sb00010100, 8'sb00010010, 8'sb00010001, 8'sb00001011, 8'sb00001100, 8'sb00010001, 8'sb00001011, 8'sb00001100, 8'sb00010100, 8'sb00010001, 8'sb00001010, 8'sb00001110, 8'sb00001001, 8'sb00010111, 8'sb00010000, 8'sb00001111, 8'sb00001101, 8'sb00001100, 8'sb00010000, 8'sb00010000, 8'sb00001110, 8'sb00000101, 8'sb11111111, 8'sb00000101, 8'sb00001000, 8'sb00001001, 8'sb00001110, 8'sb00010011, 8'sb00011010, 8'sb00001100, 8'sb00010000, 8'sb00010000, 8'sb00001110, 8'sb00001111, 8'sb00001110, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00000111, 8'sb00000001, 8'sb00000011, 8'sb00001001, 8'sb00001010, 8'sb00001111, 8'sb00001110, 8'sb00001101, 8'sb00001101,
    8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00010000, 8'sb00001101, 8'sb00010000, 8'sb00010001, 8'sb00001110, 8'sb00001101, 8'sb00001111, 8'sb00001110, 8'sb00010000, 8'sb00010001, 8'sb00010001, 8'sb00001110, 8'sb00001100, 8'sb00001101, 8'sb00001011, 8'sb00001111, 8'sb00001100, 8'sb00001101, 8'sb00010000, 8'sb00001111, 8'sb00010001, 8'sb00010000, 8'sb00001100, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00001001, 8'sb00000010, 8'sb00000001, 8'sb00010010, 8'sb00000111, 8'sb00001001, 8'sb00000100, 8'sb00001011, 8'sb00001101, 8'sb00001101, 8'sb00010001, 8'sb00010011, 8'sb00011101, 8'sb00011011, 8'sb00011000, 8'sb00011001, 8'sb00001101, 8'sb00011011, 8'sb00010011, 8'sb00010011, 8'sb00010101, 8'sb00000111, 8'sb00000111, 8'sb00001110, 8'sb00001110, 8'sb00010100, 8'sb00011101, 8'sb00011001, 8'sb00010111, 8'sb00011000, 8'sb00000110, 8'sb00101011, 8'sb00010001, 8'sb00011100, 8'sb00010101, 8'sb00001101, 8'sb00000111, 8'sb00001100, 8'sb00010010, 8'sb00011101, 8'sb00010011, 8'sb00000001, 8'sb00000011, 8'sb00001011, 8'sb00000110, 8'sb00111111, 8'sb00110111, 8'sb00100110, 8'sb00011101, 8'sb00001100, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00010101, 8'sb00000100, 8'sb00000011, 8'sb11111110, 8'sb11110110, 8'sb11101110, 8'sb00000101, 8'sb00001011, 8'sb00001001, 8'sb00001100, 8'sb00010011, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00001001, 8'sb00000000, 8'sb00000100, 8'sb11111110, 8'sb11111100, 8'sb11111101, 8'sb00000000, 8'sb00010011, 8'sb00100001, 8'sb00100001, 8'sb00001111, 8'sb00001111, 8'sb00001100, 8'sb00010001, 8'sb00001101, 8'sb00000011, 8'sb00001011, 8'sb00000000, 8'sb11111010, 8'sb00000110, 8'sb00001010, 8'sb00010001, 8'sb00011001, 8'sb00010111, 8'sb00001110, 8'sb00001110, 8'sb00010001, 8'sb00010110, 8'sb00001111, 8'sb00000001, 8'sb00001100, 8'sb00000111, 8'sb00000011, 8'sb00001100, 8'sb00001010, 8'sb00001100, 8'sb00001001, 8'sb00001011, 8'sb00001100, 8'sb00001101, 8'sb00001100, 8'sb00010100, 8'sb00010111, 8'sb00011001, 8'sb00011110, 8'sb00011000, 8'sb00100011, 8'sb00011000, 8'sb00001100, 8'sb00000000, 8'sb00000001, 8'sb11111111, 8'sb00001101, 8'sb00010001, 8'sb00001101, 8'sb00010000, 8'sb00011010, 8'sb00100101, 8'sb00010100, 8'sb00001110, 8'sb00001110, 8'sb00011000, 8'sb00010100, 8'sb00010000, 8'sb11111110, 8'sb00000011, 8'sb00001011, 8'sb00001101, 8'sb00001100, 8'sb00001110, 8'sb00010010, 8'sb00011000, 8'sb00010100, 8'sb00010010, 8'sb00010000, 8'sb00000110, 8'sb00001011, 8'sb00000111, 8'sb00000001, 8'sb00001000, 8'sb00010000, 8'sb00001110, 8'sb00001110, 8'sb00010001, 8'sb00001100, 8'sb00001100, 8'sb00001110, 8'sb00001100, 8'sb00001101, 8'sb00010110, 8'sb00010100, 8'sb00010110, 8'sb00001110, 8'sb00010000, 8'sb00010000, 8'sb00001110,
    8'sb00010011, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00001111, 8'sb00010011, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010100, 8'sb00010100, 8'sb00010001, 8'sb00001001, 8'sb00001010, 8'sb00001000, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00010011, 8'sb00010001, 8'sb00001111, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00001110, 8'sb00001101, 8'sb00000100, 8'sb00000111, 8'sb00001110, 8'sb00001100, 8'sb00010011, 8'sb00010010, 8'sb00010010, 8'sb00001110, 8'sb00010010, 8'sb00010010, 8'sb00010101, 8'sb00011011, 8'sb00010011, 8'sb00001100, 8'sb00000110, 8'sb00010011, 8'sb00010000, 8'sb00001110, 8'sb00010101, 8'sb00010011, 8'sb00010001, 8'sb00010010, 8'sb00010001, 8'sb00010000, 8'sb00010111, 8'sb00100000, 8'sb00011111, 8'sb00100000, 8'sb00010101, 8'sb00010101, 8'sb00010010, 8'sb00010010, 8'sb00010101, 8'sb00010010, 8'sb00010000, 8'sb00010001, 8'sb00001010, 8'sb00001111, 8'sb00010010, 8'sb00001100, 8'sb00010011, 8'sb00001111, 8'sb00001000, 8'sb00000101, 8'sb11111100, 8'sb11111110, 8'sb00010011, 8'sb00010100, 8'sb00010011, 8'sb00001111, 8'sb11111101, 8'sb11110001, 8'sb11101110, 8'sb11100100, 8'sb11100010, 8'sb11110101, 8'sb11111010, 8'sb11110111, 8'sb11111100, 8'sb00000000, 8'sb00001110, 8'sb00010010, 8'sb00001111, 8'sb00010000, 8'sb11110111, 8'sb11100001, 8'sb11110110, 8'sb00000011, 8'sb00010001, 8'sb00001010, 8'sb00000101, 8'sb00000111, 8'sb00010000, 8'sb00000111, 8'sb00010011, 8'sb00011001, 8'sb00010011, 8'sb00001011, 8'sb00000010, 8'sb00010000, 8'sb00011010, 8'sb00010011, 8'sb00011001, 8'sb00010101, 8'sb00001011, 8'sb00000011, 8'sb00010100, 8'sb00001110, 8'sb00011010, 8'sb00011000, 8'sb00010011, 8'sb00001101, 8'sb00010000, 8'sb00010100, 8'sb00011011, 8'sb00010101, 8'sb00011000, 8'sb00011011, 8'sb00001111, 8'sb00000111, 8'sb00000010, 8'sb00001000, 8'sb00011100, 8'sb00010101, 8'sb00001111, 8'sb00010001, 8'sb00010000, 8'sb00001100, 8'sb00010010, 8'sb00010100, 8'sb00010101, 8'sb00010110, 8'sb00001110, 8'sb00001111, 8'sb00000100, 8'sb00010100, 8'sb00011010, 8'sb00010011, 8'sb00010010, 8'sb00001111, 8'sb00001100, 8'sb00010010, 8'sb00010010, 8'sb00010010, 8'sb00010010, 8'sb00010100, 8'sb00001010, 8'sb00010001, 8'sb00010111, 8'sb00011011, 8'sb00010011, 8'sb00010000, 8'sb00010011, 8'sb00001111, 8'sb00001100, 8'sb00001000, 8'sb00001001, 8'sb00001100, 8'sb00001000, 8'sb00001100, 8'sb00010001, 8'sb00010100, 8'sb00010001, 8'sb00010001, 8'sb00010001, 8'sb00010001, 8'sb00001111, 8'sb00010010, 8'sb00010011, 8'sb00010001, 8'sb00010001, 8'sb00010110, 8'sb00010000, 8'sb00010110, 8'sb00010011, 8'sb00010000, 8'sb00010000, 8'sb00010000, 8'sb00010011, 8'sb00001111,
    8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00010010, 8'sb00001111, 8'sb00010001, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00010001, 8'sb00010001, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00001101, 8'sb00001110, 8'sb00001111, 8'sb00010001, 8'sb00010000, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00010100, 8'sb00010011, 8'sb00000110, 8'sb11111100, 8'sb11110100, 8'sb11110001, 8'sb11111001, 8'sb00000011, 8'sb00001011, 8'sb00010001, 8'sb00010000, 8'sb00001110, 8'sb00010100, 8'sb00011000, 8'sb00010101, 8'sb00011011, 8'sb00010001, 8'sb00011111, 8'sb00010001, 8'sb00010100, 8'sb00001100, 8'sb00001101, 8'sb00000101, 8'sb00001100, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00010100, 8'sb00010010, 8'sb00010100, 8'sb00011001, 8'sb00011011, 8'sb00010101, 8'sb00010010, 8'sb00011000, 8'sb00010001, 8'sb00011000, 8'sb00001010, 8'sb00010001, 8'sb00001111, 8'sb00011001, 8'sb00010001, 8'sb00001111, 8'sb00010010, 8'sb00010100, 8'sb00001111, 8'sb00010100, 8'sb00010101, 8'sb00011101, 8'sb00100011, 8'sb00010001, 8'sb00001001, 8'sb00010001, 8'sb00010011, 8'sb00010100, 8'sb00010000, 8'sb00010001, 8'sb00000101, 8'sb00001011, 8'sb00001101, 8'sb00100110, 8'sb00100000, 8'sb00010011, 8'sb00001101, 8'sb00001010, 8'sb00001010, 8'sb00010010, 8'sb00001111, 8'sb00010011, 8'sb00001001, 8'sb00000111, 8'sb00001010, 8'sb00001010, 8'sb00001110, 8'sb00010111, 8'sb00010110, 8'sb00011011, 8'sb00010101, 8'sb00001011, 8'sb00010000, 8'sb00010001, 8'sb00010000, 8'sb00010100, 8'sb00010001, 8'sb00001100, 8'sb00010000, 8'sb00001001, 8'sb00001000, 8'sb00001010, 8'sb00010100, 8'sb00010001, 8'sb00011000, 8'sb00010011, 8'sb00001110, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00001101, 8'sb11110011, 8'sb11110110, 8'sb11111010, 8'sb11111000, 8'sb00000010, 8'sb00000100, 8'sb00000110, 8'sb00010000, 8'sb00001000, 8'sb00001011, 8'sb00001110, 8'sb00010001, 8'sb00010011, 8'sb00000101, 8'sb11110011, 8'sb11111001, 8'sb11111010, 8'sb11111011, 8'sb11111101, 8'sb11111111, 8'sb00000100, 8'sb00001000, 8'sb11111110, 8'sb00001100, 8'sb00010010, 8'sb00010010, 8'sb00010011, 8'sb00010100, 8'sb00010010, 8'sb00001000, 8'sb00000111, 8'sb11111101, 8'sb00000010, 8'sb11111100, 8'sb11110110, 8'sb11111010, 8'sb00000010, 8'sb00001101, 8'sb00001110, 8'sb00010000, 8'sb00010001, 8'sb00011111, 8'sb00100101, 8'sb00010111, 8'sb00011010, 8'sb00011000, 8'sb00010000, 8'sb00010000, 8'sb00000100, 8'sb00001101, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00010001, 8'sb00010010, 8'sb00001111, 8'sb00010010, 8'sb00010010, 8'sb00010100, 8'sb00011000, 8'sb00011000, 8'sb00010110, 8'sb00010010, 8'sb00010010, 8'sb00001110, 8'sb00010001,
    8'sb00001010, 8'sb00001100, 8'sb00001101, 8'sb00001000, 8'sb00001010, 8'sb00001001, 8'sb00001011, 8'sb00001011, 8'sb00001010, 8'sb00001101, 8'sb00001100, 8'sb00001010, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00001000, 8'sb00001011, 8'sb00001000, 8'sb00001111, 8'sb00010101, 8'sb00011010, 8'sb00010011, 8'sb00010111, 8'sb00010001, 8'sb00001010, 8'sb00001110, 8'sb00001011, 8'sb00001100, 8'sb00001001, 8'sb00001010, 8'sb00000111, 8'sb00000111, 8'sb00010011, 8'sb00010001, 8'sb00000111, 8'sb00000100, 8'sb00001001, 8'sb00000011, 8'sb00001001, 8'sb00001111, 8'sb00001100, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00000101, 8'sb00010000, 8'sb00001110, 8'sb00001000, 8'sb00001111, 8'sb00001001, 8'sb00001001, 8'sb00001101, 8'sb00000100, 8'sb00001001, 8'sb00000111, 8'sb00001001, 8'sb00001010, 8'sb00001101, 8'sb00001101, 8'sb00010001, 8'sb00001001, 8'sb00010001, 8'sb00011001, 8'sb00011010, 8'sb00011010, 8'sb00001101, 8'sb00001100, 8'sb00001001, 8'sb11111101, 8'sb00001001, 8'sb00001100, 8'sb00010001, 8'sb00011111, 8'sb00011001, 8'sb00001001, 8'sb00001011, 8'sb11111111, 8'sb11111010, 8'sb00001011, 8'sb00001100, 8'sb00010011, 8'sb00011001, 8'sb00001101, 8'sb00001100, 8'sb00001001, 8'sb00010100, 8'sb00100100, 8'sb00100000, 8'sb00001000, 8'sb00001000, 8'sb11111010, 8'sb11101100, 8'sb11111110, 8'sb00000101, 8'sb00011111, 8'sb00101110, 8'sb00011100, 8'sb00001001, 8'sb00001101, 8'sb00001101, 8'sb00011111, 8'sb00110111, 8'sb00101100, 8'sb00010010, 8'sb11101111, 8'sb00000001, 8'sb00011101, 8'sb00100010, 8'sb00011011, 8'sb00010111, 8'sb00010011, 8'sb00001010, 8'sb00001010, 8'sb00001010, 8'sb00010011, 8'sb00100010, 8'sb00111111, 8'sb00111010, 8'sb00001111, 8'sb00011100, 8'sb00011101, 8'sb00010010, 8'sb00001110, 8'sb00000101, 8'sb00010010, 8'sb00001101, 8'sb00001100, 8'sb00000011, 8'sb00000101, 8'sb11111111, 8'sb00000111, 8'sb00101001, 8'sb00110010, 8'sb00010111, 8'sb00001000, 8'sb00010010, 8'sb00000110, 8'sb00001101, 8'sb00010110, 8'sb00001011, 8'sb00001010, 8'sb00001001, 8'sb00000111, 8'sb00000110, 8'sb00000010, 8'sb00001010, 8'sb00010100, 8'sb00011001, 8'sb00010010, 8'sb00001010, 8'sb00001101, 8'sb00011101, 8'sb00010100, 8'sb00001010, 8'sb00001010, 8'sb00001011, 8'sb00000111, 8'sb00001111, 8'sb00010010, 8'sb00001101, 8'sb00001011, 8'sb00000110, 8'sb00000101, 8'sb00010101, 8'sb00011010, 8'sb00011011, 8'sb00010000, 8'sb00001100, 8'sb00001001, 8'sb00001011, 8'sb00001011, 8'sb00000110, 8'sb00000011, 8'sb00000111, 8'sb00001011, 8'sb00010010, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00001100, 8'sb00001001, 8'sb00001100, 8'sb00001010, 8'sb00001010, 8'sb00001001, 8'sb00001011, 8'sb00001010, 8'sb00001101, 8'sb00010011, 8'sb00010010, 8'sb00001101, 8'sb00001111, 8'sb00001101, 8'sb00001100, 8'sb00001000, 8'sb00001100,
    8'sb00001101, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00001111, 8'sb00001110, 8'sb00010001, 8'sb00001111, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00001110, 8'sb00000100, 8'sb11111111, 8'sb00000001, 8'sb00000100, 8'sb00000011, 8'sb00000111, 8'sb00000111, 8'sb00001010, 8'sb00001110, 8'sb00010000, 8'sb00001110, 8'sb00010010, 8'sb00010011, 8'sb00010100, 8'sb00001101, 8'sb00001110, 8'sb00010111, 8'sb00010110, 8'sb00001100, 8'sb00001010, 8'sb00001001, 8'sb00001100, 8'sb00010001, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00010110, 8'sb00010000, 8'sb00010101, 8'sb00010100, 8'sb00001110, 8'sb00001000, 8'sb00000100, 8'sb11111110, 8'sb00001001, 8'sb00010101, 8'sb00010001, 8'sb00001110, 8'sb00010001, 8'sb00001110, 8'sb00011000, 8'sb00010111, 8'sb00001111, 8'sb00001100, 8'sb00001110, 8'sb00001100, 8'sb00010000, 8'sb00100000, 8'sb00011001, 8'sb00100100, 8'sb00011011, 8'sb00010001, 8'sb00001110, 8'sb00010001, 8'sb00010001, 8'sb00010001, 8'sb00010000, 8'sb00011100, 8'sb00011100, 8'sb00110000, 8'sb00100101, 8'sb00011010, 8'sb00011011, 8'sb00010100, 8'sb00011000, 8'sb00010000, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00001100, 8'sb00010111, 8'sb00010101, 8'sb00011100, 8'sb00011110, 8'sb00011010, 8'sb00010011, 8'sb00010011, 8'sb00000000, 8'sb00010000, 8'sb00010100, 8'sb00010001, 8'sb00010001, 8'sb00001100, 8'sb11111000, 8'sb00001011, 8'sb00010001, 8'sb00010101, 8'sb00011111, 8'sb00101000, 8'sb00010011, 8'sb00000011, 8'sb00000110, 8'sb00001001, 8'sb00010000, 8'sb00001111, 8'sb00011000, 8'sb00010100, 8'sb00000100, 8'sb00000010, 8'sb11111100, 8'sb00100001, 8'sb00101101, 8'sb00010000, 8'sb11111010, 8'sb00000101, 8'sb00010101, 8'sb00001110, 8'sb00001110, 8'sb00001110, 8'sb00011000, 8'sb00011000, 8'sb00010001, 8'sb00000110, 8'sb00000010, 8'sb00000110, 8'sb11111001, 8'sb11101110, 8'sb11111110, 8'sb00000001, 8'sb00001000, 8'sb00001000, 8'sb00001101, 8'sb00001101, 8'sb00010010, 8'sb00001101, 8'sb00010000, 8'sb00000111, 8'sb00000110, 8'sb00000000, 8'sb00000011, 8'sb00001001, 8'sb00000110, 8'sb00000010, 8'sb00000010, 8'sb00001000, 8'sb00001110, 8'sb00010010, 8'sb00010010, 8'sb00001100, 8'sb00010000, 8'sb00001010, 8'sb00000110, 8'sb00001111, 8'sb00010011, 8'sb00010100, 8'sb00011100, 8'sb00010101, 8'sb00010010, 8'sb00001111, 8'sb00010000, 8'sb00001111, 8'sb00010010, 8'sb00010001, 8'sb00010001, 8'sb00010101, 8'sb00010110, 8'sb00000110, 8'sb00001111, 8'sb00001110, 8'sb00010001, 8'sb00010001, 8'sb00010001, 8'sb00001111, 8'sb00001101, 8'sb00001101, 8'sb00010001, 8'sb00001101, 8'sb00001110, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00001100, 8'sb00001111, 8'sb00001100, 8'sb00001111, 8'sb00010001, 8'sb00010001, 8'sb00001101,
    8'sb00010011, 8'sb00010110, 8'sb00010101, 8'sb00010010, 8'sb00010101, 8'sb00010101, 8'sb00010011, 8'sb00010100, 8'sb00010010, 8'sb00010010, 8'sb00010011, 8'sb00010011, 8'sb00010100, 8'sb00010101, 8'sb00010110, 8'sb00010100, 8'sb00010101, 8'sb00010101, 8'sb00010001, 8'sb00001000, 8'sb00000101, 8'sb00001001, 8'sb00001010, 8'sb00001111, 8'sb00010011, 8'sb00010101, 8'sb00010010, 8'sb00010101, 8'sb00010100, 8'sb00010011, 8'sb00010011, 8'sb00010000, 8'sb00000001, 8'sb11111010, 8'sb11111101, 8'sb00000110, 8'sb00000011, 8'sb00001001, 8'sb00010010, 8'sb00011010, 8'sb00001111, 8'sb00010100, 8'sb00010011, 8'sb00010100, 8'sb00010010, 8'sb00000011, 8'sb11110111, 8'sb00000001, 8'sb00001110, 8'sb00000110, 8'sb00001000, 8'sb00010000, 8'sb00001011, 8'sb00010011, 8'sb00010101, 8'sb00010100, 8'sb00010101, 8'sb00010001, 8'sb00001110, 8'sb00000011, 8'sb11111110, 8'sb11111111, 8'sb00010110, 8'sb00011011, 8'sb00010111, 8'sb00010001, 8'sb00010000, 8'sb00001111, 8'sb00100101, 8'sb00010101, 8'sb00010010, 8'sb00010011, 8'sb00001110, 8'sb00000111, 8'sb00000111, 8'sb00001010, 8'sb00011000, 8'sb00100001, 8'sb00001011, 8'sb00000000, 8'sb00001100, 8'sb00011110, 8'sb00101101, 8'sb00010111, 8'sb00010011, 8'sb00010011, 8'sb00010110, 8'sb00010011, 8'sb00001100, 8'sb00001011, 8'sb00011000, 8'sb00010100, 8'sb00000110, 8'sb11100000, 8'sb11011101, 8'sb11101100, 8'sb00001000, 8'sb00010110, 8'sb00010101, 8'sb00010110, 8'sb00010011, 8'sb00001101, 8'sb00010010, 8'sb00001110, 8'sb00001100, 8'sb00001101, 8'sb00010000, 8'sb00001101, 8'sb11110100, 8'sb11111000, 8'sb00001101, 8'sb00010001, 8'sb00010101, 8'sb00010001, 8'sb00010010, 8'sb00001011, 8'sb00000100, 8'sb00001001, 8'sb00001101, 8'sb00010111, 8'sb00001101, 8'sb00001111, 8'sb11111001, 8'sb00000000, 8'sb00001001, 8'sb00010011, 8'sb00010110, 8'sb00010001, 8'sb00010011, 8'sb00010101, 8'sb00000111, 8'sb00001000, 8'sb00010111, 8'sb00001111, 8'sb00001100, 8'sb00010000, 8'sb11111111, 8'sb00000011, 8'sb00001101, 8'sb00010100, 8'sb00010101, 8'sb00001110, 8'sb00000100, 8'sb00001000, 8'sb00010010, 8'sb00001111, 8'sb00001001, 8'sb00001111, 8'sb00010001, 8'sb00010001, 8'sb00000100, 8'sb00001010, 8'sb00010011, 8'sb00010110, 8'sb00010101, 8'sb00010011, 8'sb00010011, 8'sb00001001, 8'sb00010011, 8'sb00001111, 8'sb00001001, 8'sb00000111, 8'sb00010101, 8'sb00011000, 8'sb00001100, 8'sb00010001, 8'sb00010010, 8'sb00010101, 8'sb00010100, 8'sb00010011, 8'sb00001110, 8'sb00001011, 8'sb00001000, 8'sb00001100, 8'sb00001010, 8'sb00000101, 8'sb00001000, 8'sb00010001, 8'sb00010000, 8'sb00010011, 8'sb00010011, 8'sb00010010, 8'sb00010100, 8'sb00010010, 8'sb00010101, 8'sb00010000, 8'sb00001110, 8'sb00010000, 8'sb00001111, 8'sb00001111, 8'sb00001100, 8'sb00010001, 8'sb00010001, 8'sb00010110, 8'sb00010110, 8'sb00010100,
    8'sb00001101, 8'sb00001011, 8'sb00001101, 8'sb00001111, 8'sb00001011, 8'sb00001111, 8'sb00001100, 8'sb00001101, 8'sb00001111, 8'sb00001101, 8'sb00001011, 8'sb00001011, 8'sb00001100, 8'sb00001011, 8'sb00001010, 8'sb00001010, 8'sb00001111, 8'sb00001110, 8'sb00010011, 8'sb00011011, 8'sb00011111, 8'sb00011111, 8'sb00011010, 8'sb00010011, 8'sb00001101, 8'sb00001101, 8'sb00001101, 8'sb00001010, 8'sb00001110, 8'sb00001101, 8'sb00001101, 8'sb00010100, 8'sb00011100, 8'sb00011011, 8'sb00011000, 8'sb00010111, 8'sb00010110, 8'sb00001101, 8'sb00000110, 8'sb00000111, 8'sb00001110, 8'sb00001111, 8'sb00001100, 8'sb00001100, 8'sb00001010, 8'sb00010000, 8'sb00010111, 8'sb00001011, 8'sb00001110, 8'sb00001001, 8'sb00000101, 8'sb00001000, 8'sb00000101, 8'sb00001000, 8'sb00010001, 8'sb00001110, 8'sb00001110, 8'sb00001001, 8'sb00000011, 8'sb00010001, 8'sb00010100, 8'sb00001011, 8'sb00000011, 8'sb00010001, 8'sb00001001, 8'sb00000111, 8'sb00010010, 8'sb00010000, 8'sb00011000, 8'sb00001101, 8'sb00001011, 8'sb00001000, 8'sb00001011, 8'sb00010001, 8'sb00000100, 8'sb00001100, 8'sb00010111, 8'sb00001100, 8'sb00000111, 8'sb00000000, 8'sb00001001, 8'sb00001010, 8'sb00010110, 8'sb00001100, 8'sb00001110, 8'sb00001011, 8'sb00000010, 8'sb11110111, 8'sb11111111, 8'sb00011000, 8'sb00010010, 8'sb11111111, 8'sb00000010, 8'sb00000111, 8'sb00000111, 8'sb00010000, 8'sb00010110, 8'sb00001011, 8'sb00001100, 8'sb00001100, 8'sb00001001, 8'sb00001000, 8'sb00001110, 8'sb00010010, 8'sb00001011, 8'sb00001110, 8'sb00000011, 8'sb00001110, 8'sb00010010, 8'sb00011010, 8'sb00100001, 8'sb00001110, 8'sb00001110, 8'sb00010001, 8'sb00011010, 8'sb00010111, 8'sb00000011, 8'sb00001001, 8'sb11111101, 8'sb00000110, 8'sb00001010, 8'sb00010011, 8'sb00001110, 8'sb00101010, 8'sb00100110, 8'sb00001110, 8'sb00001100, 8'sb00001110, 8'sb00011010, 8'sb00101001, 8'sb00101000, 8'sb00101010, 8'sb00010011, 8'sb00001100, 8'sb00010100, 8'sb00010110, 8'sb00010001, 8'sb00101100, 8'sb00011101, 8'sb00001110, 8'sb00001011, 8'sb00010000, 8'sb00011010, 8'sb00011010, 8'sb00101000, 8'sb00101111, 8'sb00100010, 8'sb00010110, 8'sb00010010, 8'sb00011000, 8'sb00010100, 8'sb00011100, 8'sb00010010, 8'sb00001110, 8'sb00001110, 8'sb00010000, 8'sb00001010, 8'sb00000001, 8'sb00001001, 8'sb00010000, 8'sb00011010, 8'sb00010110, 8'sb00010011, 8'sb00010011, 8'sb00011001, 8'sb00010000, 8'sb00001111, 8'sb00001100, 8'sb00001110, 8'sb00001101, 8'sb00000111, 8'sb00000011, 8'sb00000000, 8'sb00000010, 8'sb00000010, 8'sb00001010, 8'sb00001011, 8'sb00001011, 8'sb00000101, 8'sb00001100, 8'sb00001100, 8'sb00001011, 8'sb00001010, 8'sb00001010, 8'sb00001011, 8'sb00001101, 8'sb00001010, 8'sb00001001, 8'sb00001010, 8'sb00001000, 8'sb00001001, 8'sb00001100, 8'sb00001001, 8'sb00001100, 8'sb00001010, 8'sb00001100
    };

    localparam signed [8*30-1:0] biases_HL_param = {
    8'sb00010100, 8'sb00010011, 8'sb00010000, 8'sb00001010, 8'sb00010010, 8'sb00000011, 8'sb00000010, 8'sb00001000, 8'sb00010001, 8'sb00001101, 8'sb00001110, 8'sb00001100, 8'sb00010010, 8'sb00000100, 8'sb00011000, 8'sb00010100, 8'sb00001010, 8'sb00001111, 8'sb00010100, 8'sb00000101, 8'sb00000111, 8'sb00010010, 8'sb00001110, 8'sb00001111, 8'sb00001001, 8'sb00001001, 8'sb00010111, 8'sb00001011, 8'sb00000000, 8'sb00010010
    };

    // Instantiate the Hidden Layer
    layer #(
        .number_neuron(HL_neurons),
        .input_data_size(averaged_pixels_nr),
        .resolution(resolution)
    ) hidden_layer (
        .clk(clk), 
        .reset(reset), 
        .input_data(averaged_pixels),
        .weights(weights_HL_param),
        .biases(biases_HL_param),
        .zed(zeds_HL)
    );

    // Instantiate the Hidden Layer Sigmoid
    sigmoid_layer #(
        .number_neuron(HL_neurons)
    ) sigmoid_layer_HL (
        .zeds(zeds_HL),
        .activations(activations_HL_w)
    );

    // Instantiate dff_nbit for pixel data storage
    dff_nbit #(HL_neurons*resolution) dff_hiddel_layer (
        .clk(clk),
        .reset(reset),
        .en(1'b1),
        .di(activations_HL_w),
        .dout(activations_HL)
    );

    // Local parameters for initialized weights and biases
    localparam signed [8*10*30-1:0] weights_OL_param = {
    8'sb11000110, 8'sb10110011, 8'sb11010010, 8'sb00001001, 8'sb00101011, 8'sb11101101, 8'sb11111001, 8'sb10010111, 8'sb00011000, 8'sb11010000, 8'sb10011010, 8'sb01001111, 8'sb01000110, 8'sb00101010, 8'sb11111100, 8'sb00011101, 8'sb11110110, 8'sb00111111, 8'sb01110001, 8'sb11010100, 8'sb01011110, 8'sb11110111, 8'sb11001001, 8'sb11010010, 8'sb11011001, 8'sb00000010, 8'sb11011011, 8'sb00000101, 8'sb00010001, 8'sb11111110,
    8'sb01100111, 8'sb11111100, 8'sb11011010, 8'sb10000000, 8'sb11010110, 8'sb10011111, 8'sb11110110, 8'sb00010111, 8'sb00100110, 8'sb11001010, 8'sb11111001, 8'sb01011100, 8'sb00101011, 8'sb11110111, 8'sb00011001, 8'sb00101101, 8'sb00111111, 8'sb11010010, 8'sb11111101, 8'sb11100110, 8'sb10101000, 8'sb11101001, 8'sb01000000, 8'sb10111111, 8'sb11110110, 8'sb10110001, 8'sb11011100, 8'sb01011000, 8'sb11010101, 8'sb11011100,
    8'sb10111000, 8'sb11010010, 8'sb00001011, 8'sb11111011, 8'sb00010111, 8'sb00011010, 8'sb00111000, 8'sb01100011, 8'sb00111100, 8'sb00010011, 8'sb11111110, 8'sb11010100, 8'sb11101010, 8'sb11011010, 8'sb00010110, 8'sb11110011, 8'sb11110000, 8'sb11101110, 8'sb00001100, 8'sb00010001, 8'sb11000110, 8'sb11010101, 8'sb00000110, 8'sb01010000, 8'sb01001101, 8'sb01100010, 8'sb01010101, 8'sb11110011, 8'sb11101100, 8'sb10110110,
    8'sb00101001, 8'sb11000111, 8'sb00001111, 8'sb11001101, 8'sb11101101, 8'sb11100111, 8'sb10111010, 8'sb00110010, 8'sb10110010, 8'sb10110010, 8'sb00100011, 8'sb11101010, 8'sb00111101, 8'sb01001100, 8'sb00001011, 8'sb00001011, 8'sb11101111, 8'sb11110110, 8'sb11000111, 8'sb00110110, 8'sb00001010, 8'sb00001111, 8'sb00011101, 8'sb00000000, 8'sb11111000, 8'sb11101101, 8'sb00111110, 8'sb10111110, 8'sb00100110, 8'sb00011111,
    8'sb00011011, 8'sb00100000, 8'sb10110010, 8'sb01101100, 8'sb00111110, 8'sb00000101, 8'sb01010100, 8'sb11101011, 8'sb11001110, 8'sb11110011, 8'sb00110101, 8'sb11100010, 8'sb11010000, 8'sb11011000, 8'sb01111111, 8'sb00110001, 8'sb10001011, 8'sb00110001, 8'sb00001110, 8'sb11010000, 8'sb11101111, 8'sb11101000, 8'sb00110111, 8'sb11111001, 8'sb00101010, 8'sb11100101, 8'sb11101111, 8'sb11010001, 8'sb01110100, 8'sb11110010,
    8'sb10110000, 8'sb11010110, 8'sb00100111, 8'sb11100011, 8'sb00010110, 8'sb11100111, 8'sb00111001, 8'sb11101011, 8'sb01010001, 8'sb11100010, 8'sb01000011, 8'sb11110101, 8'sb10100111, 8'sb11111101, 8'sb11011011, 8'sb11001001, 8'sb00100101, 8'sb00010100, 8'sb10100000, 8'sb01001110, 8'sb00110011, 8'sb01010011, 8'sb00011011, 8'sb11011001, 8'sb11101100, 8'sb11101001, 8'sb11110110, 8'sb00011001, 8'sb00010100, 8'sb10111011,
    8'sb00100011, 8'sb00110000, 8'sb00110111, 8'sb01011000, 8'sb01001001, 8'sb11010001, 8'sb11001110, 8'sb10111100, 8'sb00010011, 8'sb00101001, 8'sb00001000, 8'sb11011010, 8'sb00101101, 8'sb11100010, 8'sb10011010, 8'sb11000011, 8'sb00110010, 8'sb10100110, 8'sb00011000, 8'sb00100101, 8'sb11111101, 8'sb00001111, 8'sb11010101, 8'sb00110001, 8'sb11001101, 8'sb01000001, 8'sb11001100, 8'sb00110010, 8'sb11010110, 8'sb00001010,
    8'sb11101000, 8'sb00001100, 8'sb11111110, 8'sb11101001, 8'sb11010101, 8'sb01101100, 8'sb11000010, 8'sb00100010, 8'sb11011100, 8'sb01001011, 8'sb00000001, 8'sb00100110, 8'sb11110110, 8'sb11011111, 8'sb11101100, 8'sb11010111, 8'sb00001000, 8'sb11100000, 8'sb11111011, 8'sb11010111, 8'sb00100000, 8'sb01010111, 8'sb11011001, 8'sb11101101, 8'sb01110010, 8'sb11111001, 8'sb01011010, 8'sb11101111, 8'sb11010111, 8'sb01000110,
    8'sb00010111, 8'sb00101011, 8'sb11010011, 8'sb11111011, 8'sb11111011, 8'sb01010001, 8'sb00101000, 8'sb00111011, 8'sb11000110, 8'sb00110101, 8'sb11010001, 8'sb11111011, 8'sb11111110, 8'sb01000110, 8'sb11000010, 8'sb11011011, 8'sb00000001, 8'sb11101101, 8'sb11101110, 8'sb01001000, 8'sb00111111, 8'sb11011000, 8'sb00001100, 8'sb00110000, 8'sb00001110, 8'sb11011001, 8'sb11000001, 8'sb00001111, 8'sb00111110, 8'sb11001111,
    8'sb00010100, 8'sb00000100, 8'sb00110000, 8'sb11100111, 8'sb10110011, 8'sb11101011, 8'sb11011000, 8'sb11101101, 8'sb01000100, 8'sb00000101, 8'sb00000111, 8'sb11010111, 8'sb11000110, 8'sb11110011, 8'sb00000111, 8'sb00101001, 8'sb00011110, 8'sb00110111, 8'sb00011110, 8'sb11110110, 8'sb11111100, 8'sb10111100, 8'sb11011011, 8'sb00100110, 8'sb10111010, 8'sb11100000, 8'sb01001001, 8'sb11011001, 8'sb11111000, 8'sb00100111
    };

    localparam signed [8*10-1:0] biases_OL_param = {
     8'sb11110001, 8'sb11101000, 8'sb11100111, 8'sb11100100, 8'sb11011111, 8'sb11100111, 8'sb11101110, 8'sb11101000, 8'sb11111101, 8'sb11100000
    };

    // Instantiate the Output Layer
    layer #(
        .number_neuron(OL_neurons),
        .input_data_size(HL_neurons),
        .resolution(resolution)
    ) output_layer (
        .clk(clk), 
        .reset(reset), 
        .input_data(activations_HL),
        .weights(weights_OL_param),
        .biases(biases_OL_param),
        .zed(zeds_OL)
    );

    // Instantiate the Output Layer Sigmoid
    sigmoid_layer #(
        .number_neuron(OL_neurons)
    ) sigmoid_layer_OL (
        .zeds(zeds_OL),
        .activations(activations_OL)
    );

    assign output_activations = activations_OL;

endmodule