module sigmoid(
    input wire [7:0] zed,    // 8-bit input value (unsigned)
    output reg [7:0] activation     // 8-bit activationput value (unsigned)
    );

    // Define the LUT for sigmoid values
    reg [7:0] lut [0:255];

    // Initialize the LUT with precomputed sigmoid values
    always @ * begin
        case (zed)
        -8'sd0: activation <= 8'sd0;
        -8'sd1: activation <= 8'sd0;
        -8'sd2: activation <= 8'sd0;
        -8'sd3: activation <= 8'sd0;
        -8'sd4: activation <= 8'sd0;
        -8'sd5: activation <= 8'sd0;
        -8'sd6: activation <= 8'sd0;
        -8'sd7: activation <= 8'sd0;
        -8'sd8: activation <= 8'sd0;
        -8'sd9: activation <= 8'sd0;
        -8'sd10: activation <= 8'sd0;
        -8'sd11: activation <= 8'sd0;
        -8'sd12: activation <= 8'sd0;
        -8'sd13: activation <= 8'sd0;
        -8'sd14: activation <= 8'sd0;
        -8'sd15: activation <= 8'sd0;
        -8'sd16: activation <= 8'sd0;
        -8'sd17: activation <= 8'sd0;
        -8'sd18: activation <= 8'sd1;
        -8'sd19: activation <= 8'sd1;
        -8'sd20: activation <= 8'sd1;
        -8'sd21: activation <= 8'sd1;
        -8'sd22: activation <= 8'sd1;
        -8'sd23: activation <= 8'sd1;
        -8'sd24: activation <= 8'sd1;
        -8'sd25: activation <= 8'sd1;
        -8'sd26: activation <= 8'sd1;
        -8'sd27: activation <= 8'sd1;
        -8'sd28: activation <= 8'sd1;
        -8'sd29: activation <= 8'sd1;
        -8'sd30: activation <= 8'sd1;
        -8'sd31: activation <= 8'sd1;
        -8'sd32: activation <= 8'sd2;
        -8'sd33: activation <= 8'sd2;
        -8'sd34: activation <= 8'sd2;
        -8'sd35: activation <= 8'sd2;
        -8'sd36: activation <= 8'sd2;
        -8'sd37: activation <= 8'sd2;
        -8'sd38: activation <= 8'sd2;
        -8'sd39: activation <= 8'sd2;
        -8'sd40: activation <= 8'sd3;
        -8'sd41: activation <= 8'sd3;
        -8'sd42: activation <= 8'sd3;
        -8'sd43: activation <= 8'sd3;
        -8'sd44: activation <= 8'sd3;
        -8'sd45: activation <= 8'sd3;
        -8'sd46: activation <= 8'sd4;
        -8'sd47: activation <= 8'sd4;
        -8'sd48: activation <= 8'sd4;
        -8'sd49: activation <= 8'sd4;
        -8'sd50: activation <= 8'sd5;
        -8'sd51: activation <= 8'sd5;
        -8'sd52: activation <= 8'sd5;
        -8'sd53: activation <= 8'sd5;
        -8'sd54: activation <= 8'sd6;
        -8'sd55: activation <= 8'sd6;
        -8'sd56: activation <= 8'sd6;
        -8'sd57: activation <= 8'sd7;
        -8'sd58: activation <= 8'sd7;
        -8'sd59: activation <= 8'sd7;
        -8'sd60: activation <= 8'sd8;
        -8'sd61: activation <= 8'sd8;
        -8'sd62: activation <= 8'sd9;
        -8'sd63: activation <= 8'sd9;
        -8'sd64: activation <= 8'sd9;
        -8'sd65: activation <= 8'sd10;
        -8'sd66: activation <= 8'sd10;
        -8'sd67: activation <= 8'sd11;
        -8'sd68: activation <= 8'sd12;
        -8'sd69: activation <= 8'sd12;
        -8'sd70: activation <= 8'sd13;
        -8'sd71: activation <= 8'sd13;
        -8'sd72: activation <= 8'sd14;
        -8'sd73: activation <= 8'sd15;
        -8'sd74: activation <= 8'sd16;
        -8'sd75: activation <= 8'sd16;
        -8'sd76: activation <= 8'sd17;
        -8'sd77: activation <= 8'sd18;
        -8'sd78: activation <= 8'sd19;
        -8'sd79: activation <= 8'sd20;
        -8'sd80: activation <= 8'sd21;
        -8'sd81: activation <= 8'sd22;
        -8'sd82: activation <= 8'sd23;
        -8'sd83: activation <= 8'sd24;
        -8'sd84: activation <= 8'sd25;
        -8'sd85: activation <= 8'sd26;
        -8'sd86: activation <= 8'sd27;
        -8'sd87: activation <= 8'sd29;
        -8'sd88: activation <= 8'sd30;
        -8'sd89: activation <= 8'sd31;
        -8'sd90: activation <= 8'sd33;
        -8'sd91: activation <= 8'sd34;
        -8'sd92: activation <= 8'sd36;
        -8'sd93: activation <= 8'sd37;
        -8'sd94: activation <= 8'sd39;
        -8'sd95: activation <= 8'sd41;
        -8'sd96: activation <= 8'sd42;
        -8'sd97: activation <= 8'sd44;
        -8'sd98: activation <= 8'sd46;
        -8'sd99: activation <= 8'sd48;
        -8'sd100: activation <= 8'sd50;
        -8'sd101: activation <= 8'sd52;
        -8'sd102: activation <= 8'sd54;
        -8'sd103: activation <= 8'sd56;
        -8'sd104: activation <= 8'sd59;
        -8'sd105: activation <= 8'sd61;
        -8'sd106: activation <= 8'sd63;
        -8'sd107: activation <= 8'sd66;
        -8'sd108: activation <= 8'sd68;
        -8'sd109: activation <= 8'sd71;
        -8'sd110: activation <= 8'sd73;
        -8'sd111: activation <= 8'sd76;
        -8'sd112: activation <= 8'sd79;
        -8'sd113: activation <= 8'sd81;
        -8'sd114: activation <= 8'sd84;
        -8'sd115: activation <= 8'sd87;
        -8'sd116: activation <= 8'sd90;
        -8'sd117: activation <= 8'sd93;
        -8'sd118: activation <= 8'sd96;
        -8'sd119: activation <= 8'sd99;
        -8'sd120: activation <= 8'sd102;
        -8'sd121: activation <= 8'sd105;
        -8'sd122: activation <= 8'sd108;
        -8'sd123: activation <= 8'sd111;
        -8'sd124: activation <= 8'sd114;
        -8'sd125: activation <= 8'sd117;
        -8'sd126: activation <= 8'sd121;
        -8'sd127: activation <= 8'sd124;
        8'sd128: activation <= 8'sd127;
        8'sd129: activation <= 8'sd130;
        8'sd130: activation <= 8'sd133;
        8'sd131: activation <= 8'sd137;
        8'sd132: activation <= 8'sd140;
        8'sd133: activation <= 8'sd143;
        8'sd134: activation <= 8'sd146;
        8'sd135: activation <= 8'sd149;
        8'sd136: activation <= 8'sd152;
        8'sd137: activation <= 8'sd155;
        8'sd138: activation <= 8'sd158;
        8'sd139: activation <= 8'sd161;
        8'sd140: activation <= 8'sd164;
        8'sd141: activation <= 8'sd167;
        8'sd142: activation <= 8'sd170;
        8'sd143: activation <= 8'sd173;
        8'sd144: activation <= 8'sd175;
        8'sd145: activation <= 8'sd178;
        8'sd146: activation <= 8'sd181;
        8'sd147: activation <= 8'sd183;
        8'sd148: activation <= 8'sd186;
        8'sd149: activation <= 8'sd188;
        8'sd150: activation <= 8'sd191;
        8'sd151: activation <= 8'sd193;
        8'sd152: activation <= 8'sd195;
        8'sd153: activation <= 8'sd198;
        8'sd154: activation <= 8'sd200;
        8'sd155: activation <= 8'sd202;
        8'sd156: activation <= 8'sd204;
        8'sd157: activation <= 8'sd206;
        8'sd158: activation <= 8'sd208;
        8'sd159: activation <= 8'sd210;
        8'sd160: activation <= 8'sd212;
        8'sd161: activation <= 8'sd213;
        8'sd162: activation <= 8'sd215;
        8'sd163: activation <= 8'sd217;
        8'sd164: activation <= 8'sd218;
        8'sd165: activation <= 8'sd220;
        8'sd166: activation <= 8'sd221;
        8'sd167: activation <= 8'sd223;
        8'sd168: activation <= 8'sd224;
        8'sd169: activation <= 8'sd225;
        8'sd170: activation <= 8'sd227;
        8'sd171: activation <= 8'sd228;
        8'sd172: activation <= 8'sd229;
        8'sd173: activation <= 8'sd230;
        8'sd174: activation <= 8'sd231;
        8'sd175: activation <= 8'sd232;
        8'sd176: activation <= 8'sd233;
        8'sd177: activation <= 8'sd234;
        8'sd178: activation <= 8'sd235;
        8'sd179: activation <= 8'sd236;
        8'sd180: activation <= 8'sd237;
        8'sd181: activation <= 8'sd238;
        8'sd182: activation <= 8'sd238;
        8'sd183: activation <= 8'sd239;
        8'sd184: activation <= 8'sd240;
        8'sd185: activation <= 8'sd241;
        8'sd186: activation <= 8'sd241;
        8'sd187: activation <= 8'sd242;
        8'sd188: activation <= 8'sd242;
        8'sd189: activation <= 8'sd243;
        8'sd190: activation <= 8'sd244;
        8'sd191: activation <= 8'sd244;
        8'sd192: activation <= 8'sd245;
        8'sd193: activation <= 8'sd245;
        8'sd194: activation <= 8'sd245;
        8'sd195: activation <= 8'sd246;
        8'sd196: activation <= 8'sd246;
        8'sd197: activation <= 8'sd247;
        8'sd198: activation <= 8'sd247;
        8'sd199: activation <= 8'sd247;
        8'sd200: activation <= 8'sd248;
        8'sd201: activation <= 8'sd248;
        8'sd202: activation <= 8'sd248;
        8'sd203: activation <= 8'sd249;
        8'sd204: activation <= 8'sd249;
        8'sd205: activation <= 8'sd249;
        8'sd206: activation <= 8'sd249;
        8'sd207: activation <= 8'sd250;
        8'sd208: activation <= 8'sd250;
        8'sd209: activation <= 8'sd250;
        8'sd210: activation <= 8'sd250;
        8'sd211: activation <= 8'sd251;
        8'sd212: activation <= 8'sd251;
        8'sd213: activation <= 8'sd251;
        8'sd214: activation <= 8'sd251;
        8'sd215: activation <= 8'sd251;
        8'sd216: activation <= 8'sd251;
        8'sd217: activation <= 8'sd252;
        8'sd218: activation <= 8'sd252;
        8'sd219: activation <= 8'sd252;
        8'sd220: activation <= 8'sd252;
        8'sd221: activation <= 8'sd252;
        8'sd222: activation <= 8'sd252;
        8'sd223: activation <= 8'sd252;
        8'sd224: activation <= 8'sd252;
        8'sd225: activation <= 8'sd253;
        8'sd226: activation <= 8'sd253;
        8'sd227: activation <= 8'sd253;
        8'sd228: activation <= 8'sd253;
        8'sd229: activation <= 8'sd253;
        8'sd230: activation <= 8'sd253;
        8'sd231: activation <= 8'sd253;
        8'sd232: activation <= 8'sd253;
        8'sd233: activation <= 8'sd253;
        8'sd234: activation <= 8'sd253;
        8'sd235: activation <= 8'sd253;
        8'sd236: activation <= 8'sd253;
        8'sd237: activation <= 8'sd253;
        8'sd238: activation <= 8'sd253;
        8'sd239: activation <= 8'sd254;
        8'sd240: activation <= 8'sd254;
        8'sd241: activation <= 8'sd254;
        8'sd242: activation <= 8'sd254;
        8'sd243: activation <= 8'sd254;
        8'sd244: activation <= 8'sd254;
        8'sd245: activation <= 8'sd254;
        8'sd246: activation <= 8'sd254;
        8'sd247: activation <= 8'sd254;
        8'sd248: activation <= 8'sd254;
        8'sd249: activation <= 8'sd254;
        8'sd250: activation <= 8'sd254;
        8'sd251: activation <= 8'sd254;
        8'sd252: activation <= 8'sd254;
        8'sd253: activation <= 8'sd254;
        8'sd254: activation <= 8'sd254;
        8'sd255: activation <= 8'sd254;
        endcase
    end

endmodule